module mojibake

const jis_x_0213_doublebyte_0x94 = {
	0x40: [`\u5982`].string() // U+5982 <cjk>
	0x41: [`\u5C3F`].string() // U+5C3F <cjk>
	0x42: [`\u97EE`].string() // U+97EE <cjk>
	0x43: [`\u4EFB`].string() // U+4EFB <cjk>
	0x44: [`\u598A`].string() // U+598A <cjk>
	0x45: [`\u5FCD`].string() // U+5FCD <cjk>
	0x46: [`\u8A8D`].string() // U+8A8D <cjk>
	0x47: [`\u6FE1`].string() // U+6FE1 <cjk>
	0x48: [`\u79B0`].string() // U+79B0 <cjk>
	0x49: [`\u7962`].string() // U+7962 <cjk>
	0x4A: [`\u5BE7`].string() // U+5BE7 <cjk>
	0x4B: [`\u8471`].string() // U+8471 <cjk>
	0x4C: [`\u732B`].string() // U+732B <cjk>
	0x4D: [`\u71B1`].string() // U+71B1 <cjk>
	0x4E: [`\u5E74`].string() // U+5E74 <cjk>
	0x4F: [`\u5FF5`].string() // U+5FF5 <cjk>
	0x50: [`\u637B`].string() // U+637B <cjk>
	0x51: [`\u649A`].string() // U+649A <cjk>
	0x52: [`\u71C3`].string() // U+71C3 <cjk>
	0x53: [`\u7C98`].string() // U+7C98 <cjk>
	0x54: [`\u4E43`].string() // U+4E43 <cjk>
	0x55: [`\u5EFC`].string() // U+5EFC <cjk>
	0x56: [`\u4E4B`].string() // U+4E4B <cjk>
	0x57: [`\u57DC`].string() // U+57DC <cjk>
	0x58: [`\u56A2`].string() // U+56A2 <cjk>
	0x59: [`\u60A9`].string() // U+60A9 <cjk>
	0x5A: [`\u6FC3`].string() // U+6FC3 <cjk>
	0x5B: [`\u7D0D`].string() // U+7D0D <cjk>
	0x5C: [`\u80FD`].string() // U+80FD <cjk>
	0x5D: [`\u8133`].string() // U+8133 <cjk>
	0x5E: [`\u81BF`].string() // U+81BF <cjk>
	0x5F: [`\u8FB2`].string() // U+8FB2 <cjk>
	0x60: [`\u8997`].string() // U+8997 <cjk>
	0x61: [`\u86A4`].string() // U+86A4 <cjk>
	0x62: [`\u5DF4`].string() // U+5DF4 <cjk>
	0x63: [`\u628A`].string() // U+628A <cjk>
	0x64: [`\u64AD`].string() // U+64AD <cjk>
	0x65: [`\u8987`].string() // U+8987 <cjk>
	0x66: [`\u6777`].string() // U+6777 <cjk>
	0x67: [`\u6CE2`].string() // U+6CE2 <cjk>
	0x68: [`\u6D3E`].string() // U+6D3E <cjk>
	0x69: [`\u7436`].string() // U+7436 <cjk>
	0x6A: [`\u7834`].string() // U+7834 <cjk>
	0x6B: [`\u5A46`].string() // U+5A46 <cjk>
	0x6C: [`\u7F75`].string() // U+7F75 <cjk>
	0x6D: [`\u82AD`].string() // U+82AD <cjk>
	0x6E: [`\u99AC`].string() // U+99AC <cjk>
	0x6F: [`\u4FF3`].string() // U+4FF3 <cjk>
	0x70: [`\u5EC3`].string() // U+5EC3 <cjk>
	0x71: [`\u62DD`].string() // U+62DD <cjk>
	0x72: [`\u6392`].string() // U+6392 <cjk>
	0x73: [`\u6557`].string() // U+6557 <cjk>
	0x74: [`\u676F`].string() // U+676F <cjk>
	0x75: [`\u76C3`].string() // U+76C3 <cjk>
	0x76: [`\u724C`].string() // U+724C <cjk>
	0x77: [`\u80CC`].string() // U+80CC <cjk>
	0x78: [`\u80BA`].string() // U+80BA <cjk>
	0x79: [`\u8F29`].string() // U+8F29 <cjk>
	0x7A: [`\u914D`].string() // U+914D <cjk>
	0x7B: [`\u500D`].string() // U+500D <cjk>
	0x7C: [`\u57F9`].string() // U+57F9 <cjk>
	0x7D: [`\u5A92`].string() // U+5A92 <cjk>
	0x7E: [`\u6885`].string() // U+6885 <cjk>
	0x80: [`\u6973`].string() // U+6973 <cjk>
	0x81: [`\u7164`].string() // U+7164 <cjk>
	0x82: [`\u72FD`].string() // U+72FD <cjk>
	0x83: [`\u8CB7`].string() // U+8CB7 <cjk>
	0x84: [`\u58F2`].string() // U+58F2 <cjk>
	0x85: [`\u8CE0`].string() // U+8CE0 <cjk>
	0x86: [`\u966A`].string() // U+966A <cjk>
	0x87: [`\u9019`].string() // U+9019 <cjk>
	0x88: [`\u877F`].string() // U+877F <cjk>
	0x89: [`\u79E4`].string() // U+79E4 <cjk>
	0x8A: [`\u77E7`].string() // U+77E7 <cjk>
	0x8B: [`\u8429`].string() // U+8429 <cjk>
	0x8C: [`\u4F2F`].string() // U+4F2F <cjk>
	0x8D: [`\u5265`].string() // U+5265 <cjk>
	0x8E: [`\u535A`].string() // U+535A <cjk>
	0x8F: [`\u62CD`].string() // U+62CD <cjk>
	0x90: [`\u67CF`].string() // U+67CF <cjk>
	0x91: [`\u6CCA`].string() // U+6CCA <cjk>
	0x92: [`\u767D`].string() // U+767D <cjk>
	0x93: [`\u7B94`].string() // U+7B94 <cjk>
	0x94: [`\u7C95`].string() // U+7C95 <cjk>
	0x95: [`\u8236`].string() // U+8236 <cjk>
	0x96: [`\u8584`].string() // U+8584 <cjk>
	0x97: [`\u8FEB`].string() // U+8FEB <cjk>
	0x98: [`\u66DD`].string() // U+66DD <cjk>
	0x99: [`\u6F20`].string() // U+6F20 <cjk>
	0x9A: [`\u7206`].string() // U+7206 <cjk>
	0x9B: [`\u7E1B`].string() // U+7E1B <cjk>
	0x9C: [`\u83AB`].string() // U+83AB <cjk>
	0x9D: [`\u99C1`].string() // U+99C1 <cjk>
	0x9E: [`\u9EA6`].string() // U+9EA6 <cjk>
	0x9F: [`\u51FD`].string() // U+51FD <cjk>
	0xA0: [`\u7BB1`].string() // U+7BB1 <cjk>
	0xA1: [`\u7872`].string() // U+7872 <cjk>
	0xA2: [`\u7BB8`].string() // U+7BB8 <cjk>
	0xA3: [`\u8087`].string() // U+8087 <cjk>
	0xA4: [`\u7B48`].string() // U+7B48 <cjk>
	0xA5: [`\u6AE8`].string() // U+6AE8 <cjk>
	0xA6: [`\u5E61`].string() // U+5E61 <cjk>
	0xA7: [`\u808C`].string() // U+808C <cjk>
	0xA8: [`\u7551`].string() // U+7551 <cjk>
	0xA9: [`\u7560`].string() // U+7560 <cjk>
	0xAA: [`\u516B`].string() // U+516B <cjk>
	0xAB: [`\u9262`].string() // U+9262 <cjk>
	0xAC: [`\u6E8C`].string() // U+6E8C <cjk>
	0xAD: [`\u767A`].string() // U+767A <cjk>
	0xAE: [`\u9197`].string() // U+9197 <cjk>
	0xAF: [`\u9AEA`].string() // U+9AEA <cjk>
	0xB0: [`\u4F10`].string() // U+4F10 <cjk>
	0xB1: [`\u7F70`].string() // U+7F70 <cjk>
	0xB2: [`\u629C`].string() // U+629C <cjk>
	0xB3: [`\u7B4F`].string() // U+7B4F <cjk>
	0xB4: [`\u95A5`].string() // U+95A5 <cjk>
	0xB5: [`\u9CE9`].string() // U+9CE9 <cjk>
	0xB6: [`\u567A`].string() // U+567A <cjk>
	0xB7: [`\u5859`].string() // U+5859 <cjk>
	0xB8: [`\u86E4`].string() // U+86E4 <cjk>
	0xB9: [`\u96BC`].string() // U+96BC <cjk>
	0xBA: [`\u4F34`].string() // U+4F34 <cjk>
	0xBB: [`\u5224`].string() // U+5224 <cjk>
	0xBC: [`\u534A`].string() // U+534A <cjk>
	0xBD: [`\u53CD`].string() // U+53CD <cjk>
	0xBE: [`\u53DB`].string() // U+53DB <cjk>
	0xBF: [`\u5E06`].string() // U+5E06 <cjk>
	0xC0: [`\u642C`].string() // U+642C <cjk>
	0xC1: [`\u6591`].string() // U+6591 <cjk>
	0xC2: [`\u677F`].string() // U+677F <cjk>
	0xC3: [`\u6C3E`].string() // U+6C3E <cjk>
	0xC4: [`\u6C4E`].string() // U+6C4E <cjk>
	0xC5: [`\u7248`].string() // U+7248 <cjk>
	0xC6: [`\u72AF`].string() // U+72AF <cjk>
	0xC7: [`\u73ED`].string() // U+73ED <cjk>
	0xC8: [`\u7554`].string() // U+7554 <cjk>
	0xC9: [`\u7E41`].string() // U+7E41 <cjk>
	0xCA: [`\u822C`].string() // U+822C <cjk>
	0xCB: [`\u85E9`].string() // U+85E9 <cjk>
	0xCC: [`\u8CA9`].string() // U+8CA9 <cjk>
	0xCD: [`\u7BC4`].string() // U+7BC4 <cjk>
	0xCE: [`\u91C6`].string() // U+91C6 <cjk>
	0xCF: [`\u7169`].string() // U+7169 <cjk>
	0xD0: [`\u9812`].string() // U+9812 <cjk>
	0xD1: [`\u98EF`].string() // U+98EF <cjk>
	0xD2: [`\u633D`].string() // U+633D <cjk>
	0xD3: [`\u6669`].string() // U+6669 <cjk>
	0xD4: [`\u756A`].string() // U+756A <cjk>
	0xD5: [`\u76E4`].string() // U+76E4 <cjk>
	0xD6: [`\u78D0`].string() // U+78D0 <cjk>
	0xD7: [`\u8543`].string() // U+8543 <cjk>
	0xD8: [`\u86EE`].string() // U+86EE <cjk>
	0xD9: [`\u532A`].string() // U+532A <cjk>
	0xDA: [`\u5351`].string() // U+5351 <cjk>
	0xDB: [`\u5426`].string() // U+5426 <cjk>
	0xDC: [`\u5983`].string() // U+5983 <cjk>
	0xDD: [`\u5E87`].string() // U+5E87 <cjk>
	0xDE: [`\u5F7C`].string() // U+5F7C <cjk>
	0xDF: [`\u60B2`].string() // U+60B2 <cjk>
	0xE0: [`\u6249`].string() // U+6249 <cjk>
	0xE1: [`\u6279`].string() // U+6279 <cjk>
	0xE2: [`\u62AB`].string() // U+62AB <cjk>
	0xE3: [`\u6590`].string() // U+6590 <cjk>
	0xE4: [`\u6BD4`].string() // U+6BD4 <cjk>
	0xE5: [`\u6CCC`].string() // U+6CCC <cjk>
	0xE6: [`\u75B2`].string() // U+75B2 <cjk>
	0xE7: [`\u76AE`].string() // U+76AE <cjk>
	0xE8: [`\u7891`].string() // U+7891 <cjk>
	0xE9: [`\u79D8`].string() // U+79D8 <cjk>
	0xEA: [`\u7DCB`].string() // U+7DCB <cjk>
	0xEB: [`\u7F77`].string() // U+7F77 <cjk>
	0xEC: [`\u80A5`].string() // U+80A5 <cjk>
	0xED: [`\u88AB`].string() // U+88AB <cjk>
	0xEE: [`\u8AB9`].string() // U+8AB9 <cjk>
	0xEF: [`\u8CBB`].string() // U+8CBB <cjk>
	0xF0: [`\u907F`].string() // U+907F <cjk>
	0xF1: [`\u975E`].string() // U+975E <cjk>
	0xF2: [`\u98DB`].string() // U+98DB <cjk>
	0xF3: [`\u6A0B`].string() // U+6A0B <cjk>
	0xF4: [`\u7C38`].string() // U+7C38 <cjk>
	0xF5: [`\u5099`].string() // U+5099 <cjk>
	0xF6: [`\u5C3E`].string() // U+5C3E <cjk>
	0xF7: [`\u5FAE`].string() // U+5FAE <cjk>
	0xF8: [`\u6787`].string() // U+6787 <cjk>
	0xF9: [`\u6BD8`].string() // U+6BD8 <cjk>
	0xFA: [`\u7435`].string() // U+7435 <cjk>
	0xFB: [`\u7709`].string() // U+7709 <cjk>
	0xFC: [`\u7F8E`].string() // U+7F8E <cjk>
}

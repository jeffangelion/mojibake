module mojibake

const jis_x_0213_singlebyte = {
	0x5C: [`\u00A5`].string() // U+00A5 YEN SIGN
	0x7E: [`\u203E`].string() // U+203E OVERLINE
	0xA1: [`\uFF61`].string() // U+FF61 HALFWIDTH IDEOGRAPHIC FULL STOP
	0xA2: [`\uFF62`].string() // U+FF62 HALFWIDTH LEFT CORNER BRACKET
	0xA3: [`\uFF63`].string() // U+FF63 HALFWIDTH RIGHT CORNER BRACKET
	0xA4: [`\uFF64`].string() // U+FF64 HALFWIDTH IDEOGRAPHIC COMMA
	0xA5: [`\uFF65`].string() // U+FF65 HALFWIDTH KATAKANA MIDDLE DOT
	0xA6: [`\uFF66`].string() // U+FF66 HALFWIDTH KATAKANA LETTER WO
	0xA7: [`\uFF67`].string() // U+FF67 HALFWIDTH KATAKANA LETTER SMALL A
	0xA8: [`\uFF68`].string() // U+FF68 HALFWIDTH KATAKANA LETTER SMALL I
	0xA9: [`\uFF69`].string() // U+FF69 HALFWIDTH KATAKANA LETTER SMALL U
	0xAA: [`\uFF6A`].string() // U+FF6A HALFWIDTH KATAKANA LETTER SMALL E
	0xAB: [`\uFF6B`].string() // U+FF6B HALFWIDTH KATAKANA LETTER SMALL O
	0xAC: [`\uFF6C`].string() // U+FF6C HALFWIDTH KATAKANA LETTER SMALL YA
	0xAD: [`\uFF6D`].string() // U+FF6D HALFWIDTH KATAKANA LETTER SMALL YU
	0xAE: [`\uFF6E`].string() // U+FF6E HALFWIDTH KATAKANA LETTER SMALL YO
	0xAF: [`\uFF6F`].string() // U+FF6F HALFWIDTH KATAKANA LETTER SMALL TU
	0xB0: [`\uFF70`].string() // U+FF70 HALFWIDTH KATAKANA-HIRAGANA PROLONGED SOUND MARK
	0xB1: [`\uFF71`].string() // U+FF71 HALFWIDTH KATAKANA LETTER A
	0xB2: [`\uFF72`].string() // U+FF72 HALFWIDTH KATAKANA LETTER I
	0xB3: [`\uFF73`].string() // U+FF73 HALFWIDTH KATAKANA LETTER U
	0xB4: [`\uFF74`].string() // U+FF74 HALFWIDTH KATAKANA LETTER E
	0xB5: [`\uFF75`].string() // U+FF75 HALFWIDTH KATAKANA LETTER O
	0xB6: [`\uFF76`].string() // U+FF76 HALFWIDTH KATAKANA LETTER KA
	0xB7: [`\uFF77`].string() // U+FF77 HALFWIDTH KATAKANA LETTER KI
	0xB8: [`\uFF78`].string() // U+FF78 HALFWIDTH KATAKANA LETTER KU
	0xB9: [`\uFF79`].string() // U+FF79 HALFWIDTH KATAKANA LETTER KE
	0xBA: [`\uFF7A`].string() // U+FF7A HALFWIDTH KATAKANA LETTER KO
	0xBB: [`\uFF7B`].string() // U+FF7B HALFWIDTH KATAKANA LETTER SA
	0xBC: [`\uFF7C`].string() // U+FF7C HALFWIDTH KATAKANA LETTER SI
	0xBD: [`\uFF7D`].string() // U+FF7D HALFWIDTH KATAKANA LETTER SU
	0xBE: [`\uFF7E`].string() // U+FF7E HALFWIDTH KATAKANA LETTER SE
	0xBF: [`\uFF7F`].string() // U+FF7F HALFWIDTH KATAKANA LETTER SO
	0xC0: [`\uFF80`].string() // U+FF80 HALFWIDTH KATAKANA LETTER TA
	0xC1: [`\uFF81`].string() // U+FF81 HALFWIDTH KATAKANA LETTER TI
	0xC2: [`\uFF82`].string() // U+FF82 HALFWIDTH KATAKANA LETTER TU
	0xC3: [`\uFF83`].string() // U+FF83 HALFWIDTH KATAKANA LETTER TE
	0xC4: [`\uFF84`].string() // U+FF84 HALFWIDTH KATAKANA LETTER TO
	0xC5: [`\uFF85`].string() // U+FF85 HALFWIDTH KATAKANA LETTER NA
	0xC6: [`\uFF86`].string() // U+FF86 HALFWIDTH KATAKANA LETTER NI
	0xC7: [`\uFF87`].string() // U+FF87 HALFWIDTH KATAKANA LETTER NU
	0xC8: [`\uFF88`].string() // U+FF88 HALFWIDTH KATAKANA LETTER NE
	0xC9: [`\uFF89`].string() // U+FF89 HALFWIDTH KATAKANA LETTER NO
	0xCA: [`\uFF8A`].string() // U+FF8A HALFWIDTH KATAKANA LETTER HA
	0xCB: [`\uFF8B`].string() // U+FF8B HALFWIDTH KATAKANA LETTER HI
	0xCC: [`\uFF8C`].string() // U+FF8C HALFWIDTH KATAKANA LETTER HU
	0xCD: [`\uFF8D`].string() // U+FF8D HALFWIDTH KATAKANA LETTER HE
	0xCE: [`\uFF8E`].string() // U+FF8E HALFWIDTH KATAKANA LETTER HO
	0xCF: [`\uFF8F`].string() // U+FF8F HALFWIDTH KATAKANA LETTER MA
	0xD0: [`\uFF90`].string() // U+FF90 HALFWIDTH KATAKANA LETTER MI
	0xD1: [`\uFF91`].string() // U+FF91 HALFWIDTH KATAKANA LETTER MU
	0xD2: [`\uFF92`].string() // U+FF92 HALFWIDTH KATAKANA LETTER ME
	0xD3: [`\uFF93`].string() // U+FF93 HALFWIDTH KATAKANA LETTER MO
	0xD4: [`\uFF94`].string() // U+FF94 HALFWIDTH KATAKANA LETTER YA
	0xD5: [`\uFF95`].string() // U+FF95 HALFWIDTH KATAKANA LETTER YU
	0xD6: [`\uFF96`].string() // U+FF96 HALFWIDTH KATAKANA LETTER YO
	0xD7: [`\uFF97`].string() // U+FF97 HALFWIDTH KATAKANA LETTER RA
	0xD8: [`\uFF98`].string() // U+FF98 HALFWIDTH KATAKANA LETTER RI
	0xD9: [`\uFF99`].string() // U+FF99 HALFWIDTH KATAKANA LETTER RU
	0xDA: [`\uFF9A`].string() // U+FF9A HALFWIDTH KATAKANA LETTER RE
	0xDB: [`\uFF9B`].string() // U+FF9B HALFWIDTH KATAKANA LETTER RO
	0xDC: [`\uFF9C`].string() // U+FF9C HALFWIDTH KATAKANA LETTER WA
	0xDD: [`\uFF9D`].string() // U+FF9D HALFWIDTH KATAKANA LETTER N
	0xDE: [`\uFF9E`].string() // U+FF9E HALFWIDTH KATAKANA VOICED SOUND MARK
	0xDF: [`\uFF9F`].string() // U+FF9F HALFWIDTH KATAKANA SEMI-VOICED SOUND MARK
}

module mojibake

const jis_x_0213_doublebyte_0xe0 = {
	0x40: [`\u6F3E`].string() // U+6F3E <cjk>
	0x41: [`\u6F13`].string() // U+6F13 <cjk>
	0x42: [`\u6EF7`].string() // U+6EF7 <cjk>
	0x43: [`\u6F86`].string() // U+6F86 <cjk>
	0x44: [`\u6F7A`].string() // U+6F7A <cjk>
	0x45: [`\u6F78`].string() // U+6F78 <cjk>
	0x46: [`\u6F81`].string() // U+6F81 <cjk>
	0x47: [`\u6F80`].string() // U+6F80 <cjk>
	0x48: [`\u6F6F`].string() // U+6F6F <cjk>
	0x49: [`\u6F5B`].string() // U+6F5B <cjk>
	0x4A: [`\u6FF3`].string() // U+6FF3 <cjk>
	0x4B: [`\u6F6D`].string() // U+6F6D <cjk>
	0x4C: [`\u6F82`].string() // U+6F82 <cjk>
	0x4D: [`\u6F7C`].string() // U+6F7C <cjk>
	0x4E: [`\u6F58`].string() // U+6F58 <cjk>
	0x4F: [`\u6F8E`].string() // U+6F8E <cjk>
	0x50: [`\u6F91`].string() // U+6F91 <cjk>
	0x51: [`\u6FC2`].string() // U+6FC2 <cjk>
	0x52: [`\u6F66`].string() // U+6F66 <cjk>
	0x53: [`\u6FB3`].string() // U+6FB3 <cjk>
	0x54: [`\u6FA3`].string() // U+6FA3 <cjk>
	0x55: [`\u6FA1`].string() // U+6FA1 <cjk>
	0x56: [`\u6FA4`].string() // U+6FA4 <cjk>
	0x57: [`\u6FB9`].string() // U+6FB9 <cjk>
	0x58: [`\u6FC6`].string() // U+6FC6 <cjk>
	0x59: [`\u6FAA`].string() // U+6FAA <cjk>
	0x5A: [`\u6FDF`].string() // U+6FDF <cjk>
	0x5B: [`\u6FD5`].string() // U+6FD5 <cjk>
	0x5C: [`\u6FEC`].string() // U+6FEC <cjk>
	0x5D: [`\u6FD4`].string() // U+6FD4 <cjk>
	0x5E: [`\u6FD8`].string() // U+6FD8 <cjk>
	0x5F: [`\u6FF1`].string() // U+6FF1 <cjk>
	0x60: [`\u6FEE`].string() // U+6FEE <cjk>
	0x61: [`\u6FDB`].string() // U+6FDB <cjk>
	0x62: [`\u7009`].string() // U+7009 <cjk>
	0x63: [`\u700B`].string() // U+700B <cjk>
	0x64: [`\u6FFA`].string() // U+6FFA <cjk>
	0x65: [`\u7011`].string() // U+7011 <cjk>
	0x66: [`\u7001`].string() // U+7001 <cjk>
	0x67: [`\u700F`].string() // U+700F <cjk>
	0x68: [`\u6FFE`].string() // U+6FFE <cjk>
	0x69: [`\u701B`].string() // U+701B <cjk>
	0x6A: [`\u701A`].string() // U+701A <cjk>
	0x6B: [`\u6F74`].string() // U+6F74 <cjk>
	0x6C: [`\u701D`].string() // U+701D <cjk>
	0x6D: [`\u7018`].string() // U+7018 <cjk>
	0x6E: [`\u701F`].string() // U+701F <cjk>
	0x6F: [`\u7030`].string() // U+7030 <cjk>
	0x70: [`\u703E`].string() // U+703E <cjk>
	0x71: [`\u7032`].string() // U+7032 <cjk>
	0x72: [`\u7051`].string() // U+7051 <cjk>
	0x73: [`\u7063`].string() // U+7063 <cjk>
	0x74: [`\u7099`].string() // U+7099 <cjk>
	0x75: [`\u7092`].string() // U+7092 <cjk>
	0x76: [`\u70AF`].string() // U+70AF <cjk>
	0x77: [`\u70F1`].string() // U+70F1 <cjk>
	0x78: [`\u70AC`].string() // U+70AC <cjk>
	0x79: [`\u70B8`].string() // U+70B8 <cjk>
	0x7A: [`\u70B3`].string() // U+70B3 <cjk>
	0x7B: [`\u70AE`].string() // U+70AE <cjk>
	0x7C: [`\u70DF`].string() // U+70DF <cjk>
	0x7D: [`\u70CB`].string() // U+70CB <cjk>
	0x7E: [`\u70DD`].string() // U+70DD <cjk>
	0x80: [`\u70D9`].string() // U+70D9 <cjk>
	0x81: [`\u7109`].string() // U+7109 <cjk>
	0x82: [`\u70FD`].string() // U+70FD <cjk>
	0x83: [`\u711C`].string() // U+711C <cjk>
	0x84: [`\u7119`].string() // U+7119 <cjk>
	0x85: [`\u7165`].string() // U+7165 <cjk>
	0x86: [`\u7155`].string() // U+7155 <cjk>
	0x87: [`\u7188`].string() // U+7188 <cjk>
	0x88: [`\u7166`].string() // U+7166 <cjk>
	0x89: [`\u7162`].string() // U+7162 <cjk>
	0x8A: [`\u714C`].string() // U+714C <cjk>
	0x8B: [`\u7156`].string() // U+7156 <cjk>
	0x8C: [`\u716C`].string() // U+716C <cjk>
	0x8D: [`\u718F`].string() // U+718F <cjk>
	0x8E: [`\u71FB`].string() // U+71FB <cjk>
	0x8F: [`\u7184`].string() // U+7184 <cjk>
	0x90: [`\u7195`].string() // U+7195 <cjk>
	0x91: [`\u71A8`].string() // U+71A8 <cjk>
	0x92: [`\u71AC`].string() // U+71AC <cjk>
	0x93: [`\u71D7`].string() // U+71D7 <cjk>
	0x94: [`\u71B9`].string() // U+71B9 <cjk>
	0x95: [`\u71BE`].string() // U+71BE <cjk>
	0x96: [`\u71D2`].string() // U+71D2 <cjk>
	0x97: [`\u71C9`].string() // U+71C9 <cjk>
	0x98: [`\u71D4`].string() // U+71D4 <cjk>
	0x99: [`\u71CE`].string() // U+71CE <cjk>
	0x9A: [`\u71E0`].string() // U+71E0 <cjk>
	0x9B: [`\u71EC`].string() // U+71EC <cjk>
	0x9C: [`\u71E7`].string() // U+71E7 <cjk>
	0x9D: [`\u71F5`].string() // U+71F5 <cjk>
	0x9E: [`\u71FC`].string() // U+71FC <cjk>
	0x9F: [`\u71F9`].string() // U+71F9 <cjk>
	0xA0: [`\u71FF`].string() // U+71FF <cjk>
	0xA1: [`\u720D`].string() // U+720D <cjk>
	0xA2: [`\u7210`].string() // U+7210 <cjk>
	0xA3: [`\u721B`].string() // U+721B <cjk>
	0xA4: [`\u7228`].string() // U+7228 <cjk>
	0xA5: [`\u722D`].string() // U+722D <cjk>
	0xA6: [`\u722C`].string() // U+722C <cjk>
	0xA7: [`\u7230`].string() // U+7230 <cjk>
	0xA8: [`\u7232`].string() // U+7232 <cjk>
	0xA9: [`\u723B`].string() // U+723B <cjk>
	0xAA: [`\u723C`].string() // U+723C <cjk>
	0xAB: [`\u723F`].string() // U+723F <cjk>
	0xAC: [`\u7240`].string() // U+7240 <cjk>
	0xAD: [`\u7246`].string() // U+7246 <cjk>
	0xAE: [`\u724B`].string() // U+724B <cjk>
	0xAF: [`\u7258`].string() // U+7258 <cjk>
	0xB0: [`\u7274`].string() // U+7274 <cjk>
	0xB1: [`\u727E`].string() // U+727E <cjk>
	0xB2: [`\u7282`].string() // U+7282 <cjk>
	0xB3: [`\u7281`].string() // U+7281 <cjk>
	0xB4: [`\u7287`].string() // U+7287 <cjk>
	0xB5: [`\u7292`].string() // U+7292 <cjk>
	0xB6: [`\u7296`].string() // U+7296 <cjk>
	0xB7: [`\u72A2`].string() // U+72A2 <cjk>
	0xB8: [`\u72A7`].string() // U+72A7 <cjk>
	0xB9: [`\u72B9`].string() // U+72B9 <cjk>
	0xBA: [`\u72B2`].string() // U+72B2 <cjk>
	0xBB: [`\u72C3`].string() // U+72C3 <cjk>
	0xBC: [`\u72C6`].string() // U+72C6 <cjk>
	0xBD: [`\u72C4`].string() // U+72C4 <cjk>
	0xBE: [`\u72CE`].string() // U+72CE <cjk>
	0xBF: [`\u72D2`].string() // U+72D2 <cjk>
	0xC0: [`\u72E2`].string() // U+72E2 <cjk>
	0xC1: [`\u72E0`].string() // U+72E0 <cjk>
	0xC2: [`\u72E1`].string() // U+72E1 <cjk>
	0xC3: [`\u72F9`].string() // U+72F9 <cjk>
	0xC4: [`\u72F7`].string() // U+72F7 <cjk>
	0xC5: [`\u500F`].string() // U+500F <cjk>
	0xC6: [`\u7317`].string() // U+7317 <cjk>
	0xC7: [`\u730A`].string() // U+730A <cjk>
	0xC8: [`\u731C`].string() // U+731C <cjk>
	0xC9: [`\u7316`].string() // U+7316 <cjk>
	0xCA: [`\u731D`].string() // U+731D <cjk>
	0xCB: [`\u7334`].string() // U+7334 <cjk>
	0xCC: [`\u732F`].string() // U+732F <cjk>
	0xCD: [`\u7329`].string() // U+7329 <cjk>
	0xCE: [`\u7325`].string() // U+7325 <cjk>
	0xCF: [`\u733E`].string() // U+733E <cjk>
	0xD0: [`\u734E`].string() // U+734E <cjk>
	0xD1: [`\u734F`].string() // U+734F <cjk>
	0xD2: [`\u9ED8`].string() // U+9ED8 <cjk>
	0xD3: [`\u7357`].string() // U+7357 <cjk>
	0xD4: [`\u736A`].string() // U+736A <cjk>
	0xD5: [`\u7368`].string() // U+7368 <cjk>
	0xD6: [`\u7370`].string() // U+7370 <cjk>
	0xD7: [`\u7378`].string() // U+7378 <cjk>
	0xD8: [`\u7375`].string() // U+7375 <cjk>
	0xD9: [`\u737B`].string() // U+737B <cjk>
	0xDA: [`\u737A`].string() // U+737A <cjk>
	0xDB: [`\u73C8`].string() // U+73C8 <cjk>
	0xDC: [`\u73B3`].string() // U+73B3 <cjk>
	0xDD: [`\u73CE`].string() // U+73CE <cjk>
	0xDE: [`\u73BB`].string() // U+73BB <cjk>
	0xDF: [`\u73C0`].string() // U+73C0 <cjk>
	0xE0: [`\u73E5`].string() // U+73E5 <cjk>
	0xE1: [`\u73EE`].string() // U+73EE <cjk>
	0xE2: [`\u73DE`].string() // U+73DE <cjk>
	0xE3: [`\u74A2`].string() // U+74A2 <cjk>
	0xE4: [`\u7405`].string() // U+7405 <cjk>
	0xE5: [`\u746F`].string() // U+746F <cjk>
	0xE6: [`\u7425`].string() // U+7425 <cjk>
	0xE7: [`\u73F8`].string() // U+73F8 <cjk>
	0xE8: [`\u7432`].string() // U+7432 <cjk>
	0xE9: [`\u743A`].string() // U+743A <cjk>
	0xEA: [`\u7455`].string() // U+7455 <cjk>
	0xEB: [`\u743F`].string() // U+743F <cjk>
	0xEC: [`\u745F`].string() // U+745F <cjk>
	0xED: [`\u7459`].string() // U+7459 <cjk>
	0xEE: [`\u7441`].string() // U+7441 <cjk>
	0xEF: [`\u745C`].string() // U+745C <cjk>
	0xF0: [`\u7469`].string() // U+7469 <cjk>
	0xF1: [`\u7470`].string() // U+7470 <cjk>
	0xF2: [`\u7463`].string() // U+7463 <cjk>
	0xF3: [`\u746A`].string() // U+746A <cjk>
	0xF4: [`\u7476`].string() // U+7476 <cjk>
	0xF5: [`\u747E`].string() // U+747E <cjk>
	0xF6: [`\u748B`].string() // U+748B <cjk>
	0xF7: [`\u749E`].string() // U+749E <cjk>
	0xF8: [`\u74A7`].string() // U+74A7 <cjk>
	0xF9: [`\u74CA`].string() // U+74CA <cjk>
	0xFA: [`\u74CF`].string() // U+74CF <cjk>
	0xFB: [`\u74D4`].string() // U+74D4 <cjk>
	0xFC: [`\u73F1`].string() // U+73F1 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x8c = {
	0x40: [`\u6398`].string() // U+6398 <cjk>
	0x41: [`\u7A9F`].string() // U+7A9F <cjk>
	0x42: [`\u6C93`].string() // U+6C93 <cjk>
	0x43: [`\u9774`].string() // U+9774 <cjk>
	0x44: [`\u8F61`].string() // U+8F61 <cjk>
	0x45: [`\u7AAA`].string() // U+7AAA <cjk>
	0x46: [`\u718A`].string() // U+718A <cjk>
	0x47: [`\u9688`].string() // U+9688 <cjk>
	0x48: [`\u7C82`].string() // U+7C82 <cjk>
	0x49: [`\u6817`].string() // U+6817 <cjk>
	0x4A: [`\u7E70`].string() // U+7E70 <cjk>
	0x4B: [`\u6851`].string() // U+6851 <cjk>
	0x4C: [`\u936C`].string() // U+936C <cjk>
	0x4D: [`\u52F2`].string() // U+52F2 <cjk>
	0x4E: [`\u541B`].string() // U+541B <cjk>
	0x4F: [`\u85AB`].string() // U+85AB <cjk>
	0x50: [`\u8A13`].string() // U+8A13 <cjk>
	0x51: [`\u7FA4`].string() // U+7FA4 <cjk>
	0x52: [`\u8ECD`].string() // U+8ECD <cjk>
	0x53: [`\u90E1`].string() // U+90E1 <cjk>
	0x54: [`\u5366`].string() // U+5366 <cjk>
	0x55: [`\u8888`].string() // U+8888 <cjk>
	0x56: [`\u7941`].string() // U+7941 <cjk>
	0x57: [`\u4FC2`].string() // U+4FC2 <cjk>
	0x58: [`\u50BE`].string() // U+50BE <cjk>
	0x59: [`\u5211`].string() // U+5211 <cjk>
	0x5A: [`\u5144`].string() // U+5144 <cjk>
	0x5B: [`\u5553`].string() // U+5553 <cjk>
	0x5C: [`\u572D`].string() // U+572D <cjk>
	0x5D: [`\u73EA`].string() // U+73EA <cjk>
	0x5E: [`\u578B`].string() // U+578B <cjk>
	0x5F: [`\u5951`].string() // U+5951 <cjk>
	0x60: [`\u5F62`].string() // U+5F62 <cjk>
	0x61: [`\u5F84`].string() // U+5F84 <cjk>
	0x62: [`\u6075`].string() // U+6075 <cjk>
	0x63: [`\u6176`].string() // U+6176 <cjk>
	0x64: [`\u6167`].string() // U+6167 <cjk>
	0x65: [`\u61A9`].string() // U+61A9 <cjk>
	0x66: [`\u63B2`].string() // U+63B2 <cjk>
	0x67: [`\u643A`].string() // U+643A <cjk>
	0x68: [`\u656C`].string() // U+656C <cjk>
	0x69: [`\u666F`].string() // U+666F <cjk>
	0x6A: [`\u6842`].string() // U+6842 <cjk>
	0x6B: [`\u6E13`].string() // U+6E13 <cjk>
	0x6C: [`\u7566`].string() // U+7566 <cjk>
	0x6D: [`\u7A3D`].string() // U+7A3D <cjk>
	0x6E: [`\u7CFB`].string() // U+7CFB <cjk>
	0x6F: [`\u7D4C`].string() // U+7D4C <cjk>
	0x70: [`\u7D99`].string() // U+7D99 <cjk>
	0x71: [`\u7E4B`].string() // U+7E4B <cjk>
	0x72: [`\u7F6B`].string() // U+7F6B <cjk>
	0x73: [`\u830E`].string() // U+830E <cjk>
	0x74: [`\u834A`].string() // U+834A <cjk>
	0x75: [`\u86CD`].string() // U+86CD <cjk>
	0x76: [`\u8A08`].string() // U+8A08 <cjk>
	0x77: [`\u8A63`].string() // U+8A63 <cjk>
	0x78: [`\u8B66`].string() // U+8B66 <cjk>
	0x79: [`\u8EFD`].string() // U+8EFD <cjk>
	0x7A: [`\u981A`].string() // U+981A <cjk>
	0x7B: [`\u9D8F`].string() // U+9D8F <cjk>
	0x7C: [`\u82B8`].string() // U+82B8 <cjk>
	0x7D: [`\u8FCE`].string() // U+8FCE <cjk>
	0x7E: [`\u9BE8`].string() // U+9BE8 <cjk>
	0x80: [`\u5287`].string() // U+5287 <cjk>
	0x81: [`\u621F`].string() // U+621F <cjk>
	0x82: [`\u6483`].string() // U+6483 <cjk>
	0x83: [`\u6FC0`].string() // U+6FC0 <cjk>
	0x84: [`\u9699`].string() // U+9699 <cjk>
	0x85: [`\u6841`].string() // U+6841 <cjk>
	0x86: [`\u5091`].string() // U+5091 <cjk>
	0x87: [`\u6B20`].string() // U+6B20 <cjk>
	0x88: [`\u6C7A`].string() // U+6C7A <cjk>
	0x89: [`\u6F54`].string() // U+6F54 <cjk>
	0x8A: [`\u7A74`].string() // U+7A74 <cjk>
	0x8B: [`\u7D50`].string() // U+7D50 <cjk>
	0x8C: [`\u8840`].string() // U+8840 <cjk>
	0x8D: [`\u8A23`].string() // U+8A23 <cjk>
	0x8E: [`\u6708`].string() // U+6708 <cjk>
	0x8F: [`\u4EF6`].string() // U+4EF6 <cjk>
	0x90: [`\u5039`].string() // U+5039 <cjk>
	0x91: [`\u5026`].string() // U+5026 <cjk>
	0x92: [`\u5065`].string() // U+5065 <cjk>
	0x93: [`\u517C`].string() // U+517C <cjk>
	0x94: [`\u5238`].string() // U+5238 <cjk>
	0x95: [`\u5263`].string() // U+5263 <cjk>
	0x96: [`\u55A7`].string() // U+55A7 <cjk>
	0x97: [`\u570F`].string() // U+570F <cjk>
	0x98: [`\u5805`].string() // U+5805 <cjk>
	0x99: [`\u5ACC`].string() // U+5ACC <cjk>
	0x9A: [`\u5EFA`].string() // U+5EFA <cjk>
	0x9B: [`\u61B2`].string() // U+61B2 <cjk>
	0x9C: [`\u61F8`].string() // U+61F8 <cjk>
	0x9D: [`\u62F3`].string() // U+62F3 <cjk>
	0x9E: [`\u6372`].string() // U+6372 <cjk>
	0x9F: [`\u691C`].string() // U+691C <cjk>
	0xA0: [`\u6A29`].string() // U+6A29 <cjk>
	0xA1: [`\u727D`].string() // U+727D <cjk>
	0xA2: [`\u72AC`].string() // U+72AC <cjk>
	0xA3: [`\u732E`].string() // U+732E <cjk>
	0xA4: [`\u7814`].string() // U+7814 <cjk>
	0xA5: [`\u786F`].string() // U+786F <cjk>
	0xA6: [`\u7D79`].string() // U+7D79 <cjk>
	0xA7: [`\u770C`].string() // U+770C <cjk>
	0xA8: [`\u80A9`].string() // U+80A9 <cjk>
	0xA9: [`\u898B`].string() // U+898B <cjk>
	0xAA: [`\u8B19`].string() // U+8B19 <cjk>
	0xAB: [`\u8CE2`].string() // U+8CE2 <cjk>
	0xAC: [`\u8ED2`].string() // U+8ED2 <cjk>
	0xAD: [`\u9063`].string() // U+9063 <cjk>
	0xAE: [`\u9375`].string() // U+9375 <cjk>
	0xAF: [`\u967A`].string() // U+967A <cjk>
	0xB0: [`\u9855`].string() // U+9855 <cjk>
	0xB1: [`\u9A13`].string() // U+9A13 <cjk>
	0xB2: [`\u9E78`].string() // U+9E78 <cjk>
	0xB3: [`\u5143`].string() // U+5143 <cjk>
	0xB4: [`\u539F`].string() // U+539F <cjk>
	0xB5: [`\u53B3`].string() // U+53B3 <cjk>
	0xB6: [`\u5E7B`].string() // U+5E7B <cjk>
	0xB7: [`\u5F26`].string() // U+5F26 <cjk>
	0xB8: [`\u6E1B`].string() // U+6E1B <cjk>
	0xB9: [`\u6E90`].string() // U+6E90 <cjk>
	0xBA: [`\u7384`].string() // U+7384 <cjk>
	0xBB: [`\u73FE`].string() // U+73FE <cjk>
	0xBC: [`\u7D43`].string() // U+7D43 <cjk>
	0xBD: [`\u8237`].string() // U+8237 <cjk>
	0xBE: [`\u8A00`].string() // U+8A00 <cjk>
	0xBF: [`\u8AFA`].string() // U+8AFA <cjk>
	0xC0: [`\u9650`].string() // U+9650 <cjk>
	0xC1: [`\u4E4E`].string() // U+4E4E <cjk>
	0xC2: [`\u500B`].string() // U+500B <cjk>
	0xC3: [`\u53E4`].string() // U+53E4 <cjk>
	0xC4: [`\u547C`].string() // U+547C <cjk>
	0xC5: [`\u56FA`].string() // U+56FA <cjk>
	0xC6: [`\u59D1`].string() // U+59D1 <cjk>
	0xC7: [`\u5B64`].string() // U+5B64 <cjk>
	0xC8: [`\u5DF1`].string() // U+5DF1 <cjk>
	0xC9: [`\u5EAB`].string() // U+5EAB <cjk>
	0xCA: [`\u5F27`].string() // U+5F27 <cjk>
	0xCB: [`\u6238`].string() // U+6238 <cjk>
	0xCC: [`\u6545`].string() // U+6545 <cjk>
	0xCD: [`\u67AF`].string() // U+67AF <cjk>
	0xCE: [`\u6E56`].string() // U+6E56 <cjk>
	0xCF: [`\u72D0`].string() // U+72D0 <cjk>
	0xD0: [`\u7CCA`].string() // U+7CCA <cjk>
	0xD1: [`\u88B4`].string() // U+88B4 <cjk>
	0xD2: [`\u80A1`].string() // U+80A1 <cjk>
	0xD3: [`\u80E1`].string() // U+80E1 <cjk>
	0xD4: [`\u83F0`].string() // U+83F0 <cjk>
	0xD5: [`\u864E`].string() // U+864E <cjk>
	0xD6: [`\u8A87`].string() // U+8A87 <cjk>
	0xD7: [`\u8DE8`].string() // U+8DE8 <cjk>
	0xD8: [`\u9237`].string() // U+9237 <cjk>
	0xD9: [`\u96C7`].string() // U+96C7 <cjk>
	0xDA: [`\u9867`].string() // U+9867 <cjk>
	0xDB: [`\u9F13`].string() // U+9F13 <cjk>
	0xDC: [`\u4E94`].string() // U+4E94 <cjk>
	0xDD: [`\u4E92`].string() // U+4E92 <cjk>
	0xDE: [`\u4F0D`].string() // U+4F0D <cjk>
	0xDF: [`\u5348`].string() // U+5348 <cjk>
	0xE0: [`\u5449`].string() // U+5449 <cjk>
	0xE1: [`\u543E`].string() // U+543E <cjk>
	0xE2: [`\u5A2F`].string() // U+5A2F <cjk>
	0xE3: [`\u5F8C`].string() // U+5F8C <cjk>
	0xE4: [`\u5FA1`].string() // U+5FA1 <cjk>
	0xE5: [`\u609F`].string() // U+609F <cjk>
	0xE6: [`\u68A7`].string() // U+68A7 <cjk>
	0xE7: [`\u6A8E`].string() // U+6A8E <cjk>
	0xE8: [`\u745A`].string() // U+745A <cjk>
	0xE9: [`\u7881`].string() // U+7881 <cjk>
	0xEA: [`\u8A9E`].string() // U+8A9E <cjk>
	0xEB: [`\u8AA4`].string() // U+8AA4 <cjk>
	0xEC: [`\u8B77`].string() // U+8B77 <cjk>
	0xED: [`\u9190`].string() // U+9190 <cjk>
	0xEE: [`\u4E5E`].string() // U+4E5E <cjk>
	0xEF: [`\u9BC9`].string() // U+9BC9 <cjk>
	0xF0: [`\u4EA4`].string() // U+4EA4 <cjk>
	0xF1: [`\u4F7C`].string() // U+4F7C <cjk>
	0xF2: [`\u4FAF`].string() // U+4FAF <cjk>
	0xF3: [`\u5019`].string() // U+5019 <cjk>
	0xF4: [`\u5016`].string() // U+5016 <cjk>
	0xF5: [`\u5149`].string() // U+5149 <cjk>
	0xF6: [`\u516C`].string() // U+516C <cjk>
	0xF7: [`\u529F`].string() // U+529F <cjk>
	0xF8: [`\u52B9`].string() // U+52B9 <cjk>
	0xF9: [`\u52FE`].string() // U+52FE <cjk>
	0xFA: [`\u539A`].string() // U+539A <cjk>
	0xFB: [`\u53E3`].string() // U+53E3 <cjk>
	0xFC: [`\u5411`].string() // U+5411 <cjk>
}

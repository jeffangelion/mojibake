module mojibake

const jis_x_0213_doublebyte_0x97 = {
	0x40: [`\u8AED`].string() // U+8AED <cjk>
	0x41: [`\u8F38`].string() // U+8F38 <cjk>
	0x42: [`\u552F`].string() // U+552F <cjk>
	0x43: [`\u4F51`].string() // U+4F51 <cjk>
	0x44: [`\u512A`].string() // U+512A <cjk>
	0x45: [`\u52C7`].string() // U+52C7 <cjk>
	0x46: [`\u53CB`].string() // U+53CB <cjk>
	0x47: [`\u5BA5`].string() // U+5BA5 <cjk>
	0x48: [`\u5E7D`].string() // U+5E7D <cjk>
	0x49: [`\u60A0`].string() // U+60A0 <cjk>
	0x4A: [`\u6182`].string() // U+6182 <cjk>
	0x4B: [`\u63D6`].string() // U+63D6 <cjk>
	0x4C: [`\u6709`].string() // U+6709 <cjk>
	0x4D: [`\u67DA`].string() // U+67DA <cjk>
	0x4E: [`\u6E67`].string() // U+6E67 <cjk>
	0x4F: [`\u6D8C`].string() // U+6D8C <cjk>
	0x50: [`\u7336`].string() // U+7336 <cjk>
	0x51: [`\u7337`].string() // U+7337 <cjk>
	0x52: [`\u7531`].string() // U+7531 <cjk>
	0x53: [`\u7950`].string() // U+7950 <cjk>
	0x54: [`\u88D5`].string() // U+88D5 <cjk>
	0x55: [`\u8A98`].string() // U+8A98 <cjk>
	0x56: [`\u904A`].string() // U+904A <cjk>
	0x57: [`\u9091`].string() // U+9091 <cjk>
	0x58: [`\u90F5`].string() // U+90F5 <cjk>
	0x59: [`\u96C4`].string() // U+96C4 <cjk>
	0x5A: [`\u878D`].string() // U+878D <cjk>
	0x5B: [`\u5915`].string() // U+5915 <cjk>
	0x5C: [`\u4E88`].string() // U+4E88 <cjk>
	0x5D: [`\u4F59`].string() // U+4F59 <cjk>
	0x5E: [`\u4E0E`].string() // U+4E0E <cjk>
	0x5F: [`\u8A89`].string() // U+8A89 <cjk>
	0x60: [`\u8F3F`].string() // U+8F3F <cjk>
	0x61: [`\u9810`].string() // U+9810 <cjk>
	0x62: [`\u50AD`].string() // U+50AD <cjk>
	0x63: [`\u5E7C`].string() // U+5E7C <cjk>
	0x64: [`\u5996`].string() // U+5996 <cjk>
	0x65: [`\u5BB9`].string() // U+5BB9 <cjk>
	0x66: [`\u5EB8`].string() // U+5EB8 <cjk>
	0x67: [`\u63DA`].string() // U+63DA <cjk>
	0x68: [`\u63FA`].string() // U+63FA <cjk>
	0x69: [`\u64C1`].string() // U+64C1 <cjk>
	0x6A: [`\u66DC`].string() // U+66DC <cjk>
	0x6B: [`\u694A`].string() // U+694A <cjk>
	0x6C: [`\u69D8`].string() // U+69D8 <cjk>
	0x6D: [`\u6D0B`].string() // U+6D0B <cjk>
	0x6E: [`\u6EB6`].string() // U+6EB6 <cjk>
	0x6F: [`\u7194`].string() // U+7194 <cjk>
	0x70: [`\u7528`].string() // U+7528 <cjk>
	0x71: [`\u7AAF`].string() // U+7AAF <cjk>
	0x72: [`\u7F8A`].string() // U+7F8A <cjk>
	0x73: [`\u8000`].string() // U+8000 <cjk>
	0x74: [`\u8449`].string() // U+8449 <cjk>
	0x75: [`\u84C9`].string() // U+84C9 <cjk>
	0x76: [`\u8981`].string() // U+8981 <cjk>
	0x77: [`\u8B21`].string() // U+8B21 <cjk>
	0x78: [`\u8E0A`].string() // U+8E0A <cjk>
	0x79: [`\u9065`].string() // U+9065 <cjk>
	0x7A: [`\u967D`].string() // U+967D <cjk>
	0x7B: [`\u990A`].string() // U+990A <cjk>
	0x7C: [`\u617E`].string() // U+617E <cjk>
	0x7D: [`\u6291`].string() // U+6291 <cjk>
	0x7E: [`\u6B32`].string() // U+6B32 <cjk>
	0x80: [`\u6C83`].string() // U+6C83 <cjk>
	0x81: [`\u6D74`].string() // U+6D74 <cjk>
	0x82: [`\u7FCC`].string() // U+7FCC <cjk>
	0x83: [`\u7FFC`].string() // U+7FFC <cjk>
	0x84: [`\u6DC0`].string() // U+6DC0 <cjk>
	0x85: [`\u7F85`].string() // U+7F85 <cjk>
	0x86: [`\u87BA`].string() // U+87BA <cjk>
	0x87: [`\u88F8`].string() // U+88F8 <cjk>
	0x88: [`\u6765`].string() // U+6765 <cjk>
	0x89: [`\u83B1`].string() // U+83B1 <cjk>
	0x8A: [`\u983C`].string() // U+983C <cjk>
	0x8B: [`\u96F7`].string() // U+96F7 <cjk>
	0x8C: [`\u6D1B`].string() // U+6D1B <cjk>
	0x8D: [`\u7D61`].string() // U+7D61 <cjk>
	0x8E: [`\u843D`].string() // U+843D <cjk>
	0x8F: [`\u916A`].string() // U+916A <cjk>
	0x90: [`\u4E71`].string() // U+4E71 <cjk>
	0x91: [`\u5375`].string() // U+5375 <cjk>
	0x92: [`\u5D50`].string() // U+5D50 <cjk>
	0x93: [`\u6B04`].string() // U+6B04 <cjk>
	0x94: [`\u6FEB`].string() // U+6FEB <cjk>
	0x95: [`\u85CD`].string() // U+85CD <cjk>
	0x96: [`\u862D`].string() // U+862D <cjk>
	0x97: [`\u89A7`].string() // U+89A7 <cjk>
	0x98: [`\u5229`].string() // U+5229 <cjk>
	0x99: [`\u540F`].string() // U+540F <cjk>
	0x9A: [`\u5C65`].string() // U+5C65 <cjk>
	0x9B: [`\u674E`].string() // U+674E <cjk>
	0x9C: [`\u68A8`].string() // U+68A8 <cjk>
	0x9D: [`\u7406`].string() // U+7406 <cjk>
	0x9E: [`\u7483`].string() // U+7483 <cjk>
	0x9F: [`\u75E2`].string() // U+75E2 <cjk>
	0xA0: [`\u88CF`].string() // U+88CF <cjk>
	0xA1: [`\u88E1`].string() // U+88E1 <cjk>
	0xA2: [`\u91CC`].string() // U+91CC <cjk>
	0xA3: [`\u96E2`].string() // U+96E2 <cjk>
	0xA4: [`\u9678`].string() // U+9678 <cjk>
	0xA5: [`\u5F8B`].string() // U+5F8B <cjk>
	0xA6: [`\u7387`].string() // U+7387 <cjk>
	0xA7: [`\u7ACB`].string() // U+7ACB <cjk>
	0xA8: [`\u844E`].string() // U+844E <cjk>
	0xA9: [`\u63A0`].string() // U+63A0 <cjk>
	0xAA: [`\u7565`].string() // U+7565 <cjk>
	0xAB: [`\u5289`].string() // U+5289 <cjk>
	0xAC: [`\u6D41`].string() // U+6D41 <cjk>
	0xAD: [`\u6E9C`].string() // U+6E9C <cjk>
	0xAE: [`\u7409`].string() // U+7409 <cjk>
	0xAF: [`\u7559`].string() // U+7559 <cjk>
	0xB0: [`\u786B`].string() // U+786B <cjk>
	0xB1: [`\u7C92`].string() // U+7C92 <cjk>
	0xB2: [`\u9686`].string() // U+9686 <cjk>
	0xB3: [`\u7ADC`].string() // U+7ADC <cjk>
	0xB4: [`\u9F8D`].string() // U+9F8D <cjk>
	0xB5: [`\u4FB6`].string() // U+4FB6 <cjk>
	0xB6: [`\u616E`].string() // U+616E <cjk>
	0xB7: [`\u65C5`].string() // U+65C5 <cjk>
	0xB8: [`\u865C`].string() // U+865C <cjk>
	0xB9: [`\u4E86`].string() // U+4E86 <cjk>
	0xBA: [`\u4EAE`].string() // U+4EAE <cjk>
	0xBB: [`\u50DA`].string() // U+50DA <cjk>
	0xBC: [`\u4E21`].string() // U+4E21 <cjk>
	0xBD: [`\u51CC`].string() // U+51CC <cjk>
	0xBE: [`\u5BEE`].string() // U+5BEE <cjk>
	0xBF: [`\u6599`].string() // U+6599 <cjk>
	0xC0: [`\u6881`].string() // U+6881 <cjk>
	0xC1: [`\u6DBC`].string() // U+6DBC <cjk>
	0xC2: [`\u731F`].string() // U+731F <cjk>
	0xC3: [`\u7642`].string() // U+7642 <cjk>
	0xC4: [`\u77AD`].string() // U+77AD <cjk>
	0xC5: [`\u7A1C`].string() // U+7A1C <cjk>
	0xC6: [`\u7CE7`].string() // U+7CE7 <cjk>
	0xC7: [`\u826F`].string() // U+826F <cjk>
	0xC8: [`\u8AD2`].string() // U+8AD2 <cjk>
	0xC9: [`\u907C`].string() // U+907C <cjk>
	0xCA: [`\u91CF`].string() // U+91CF <cjk>
	0xCB: [`\u9675`].string() // U+9675 <cjk>
	0xCC: [`\u9818`].string() // U+9818 <cjk>
	0xCD: [`\u529B`].string() // U+529B <cjk>
	0xCE: [`\u7DD1`].string() // U+7DD1 <cjk>
	0xCF: [`\u502B`].string() // U+502B <cjk>
	0xD0: [`\u5398`].string() // U+5398 <cjk>
	0xD1: [`\u6797`].string() // U+6797 <cjk>
	0xD2: [`\u6DCB`].string() // U+6DCB <cjk>
	0xD3: [`\u71D0`].string() // U+71D0 <cjk>
	0xD4: [`\u7433`].string() // U+7433 <cjk>
	0xD5: [`\u81E8`].string() // U+81E8 <cjk>
	0xD6: [`\u8F2A`].string() // U+8F2A <cjk>
	0xD7: [`\u96A3`].string() // U+96A3 <cjk>
	0xD8: [`\u9C57`].string() // U+9C57 <cjk>
	0xD9: [`\u9E9F`].string() // U+9E9F <cjk>
	0xDA: [`\u7460`].string() // U+7460 <cjk>
	0xDB: [`\u5841`].string() // U+5841 <cjk>
	0xDC: [`\u6D99`].string() // U+6D99 <cjk>
	0xDD: [`\u7D2F`].string() // U+7D2F <cjk>
	0xDE: [`\u985E`].string() // U+985E <cjk>
	0xDF: [`\u4EE4`].string() // U+4EE4 <cjk>
	0xE0: [`\u4F36`].string() // U+4F36 <cjk>
	0xE1: [`\u4F8B`].string() // U+4F8B <cjk>
	0xE2: [`\u51B7`].string() // U+51B7 <cjk>
	0xE3: [`\u52B1`].string() // U+52B1 <cjk>
	0xE4: [`\u5DBA`].string() // U+5DBA <cjk>
	0xE5: [`\u601C`].string() // U+601C <cjk>
	0xE6: [`\u73B2`].string() // U+73B2 <cjk>
	0xE7: [`\u793C`].string() // U+793C <cjk>
	0xE8: [`\u82D3`].string() // U+82D3 <cjk>
	0xE9: [`\u9234`].string() // U+9234 <cjk>
	0xEA: [`\u96B7`].string() // U+96B7 <cjk>
	0xEB: [`\u96F6`].string() // U+96F6 <cjk>
	0xEC: [`\u970A`].string() // U+970A <cjk>
	0xED: [`\u9E97`].string() // U+9E97 <cjk>
	0xEE: [`\u9F62`].string() // U+9F62 <cjk>
	0xEF: [`\u66A6`].string() // U+66A6 <cjk>
	0xF0: [`\u6B74`].string() // U+6B74 <cjk>
	0xF1: [`\u5217`].string() // U+5217 <cjk>
	0xF2: [`\u52A3`].string() // U+52A3 <cjk>
	0xF3: [`\u70C8`].string() // U+70C8 <cjk>
	0xF4: [`\u88C2`].string() // U+88C2 <cjk>
	0xF5: [`\u5EC9`].string() // U+5EC9 <cjk>
	0xF6: [`\u604B`].string() // U+604B <cjk>
	0xF7: [`\u6190`].string() // U+6190 <cjk>
	0xF8: [`\u6F23`].string() // U+6F23 <cjk>
	0xF9: [`\u7149`].string() // U+7149 <cjk>
	0xFA: [`\u7C3E`].string() // U+7C3E <cjk>
	0xFB: [`\u7DF4`].string() // U+7DF4 <cjk>
	0xFC: [`\u806F`].string() // U+806F <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xeb = {
	0x40: [`\u64C4`].string() // U+64C4 <cjk>
	0x41: [`\u64CA`].string() // U+64CA <cjk>
	0x42: [`\u64D0`].string() // U+64D0 <cjk>
	0x43: [`\u64F7`].string() // U+64F7 <cjk>
	0x44: [`\u64FB`].string() // U+64FB <cjk>
	0x45: [`\u6522`].string() // U+6522 <cjk>
	0x46: [`\u6529`].string() // U+6529 <cjk>
	0x47: [`\uFA41`].string() // U+FA41 CJK COMPATIBILITY IDEOGRAPH-FA41
	0x48: [`\u6567`].string() // U+6567 <cjk>
	0x49: [`\u659D`].string() // U+659D <cjk>
	0x4A: [`\uFA42`].string() // U+FA42 CJK COMPATIBILITY IDEOGRAPH-FA42
	0x4B: [`\u6600`].string() // U+6600 <cjk>
	0x4C: [`\u6609`].string() // U+6609 <cjk>
	0x4D: [`\u6615`].string() // U+6615 <cjk>
	0x4E: [`\u661E`].string() // U+661E <cjk>
	0x4F: [`\u663A`].string() // U+663A <cjk>
	0x50: [`\u6622`].string() // U+6622 <cjk>
	0x51: [`\u6624`].string() // U+6624 <cjk>
	0x52: [`\u662B`].string() // U+662B <cjk>
	0x53: [`\u6630`].string() // U+6630 <cjk>
	0x54: [`\u6631`].string() // U+6631 <cjk>
	0x55: [`\u6633`].string() // U+6633 <cjk>
	0x56: [`\u66FB`].string() // U+66FB <cjk>
	0x57: [`\u6648`].string() // U+6648 <cjk>
	0x58: [`\u664C`].string() // U+664C <cjk>
	0x59: utf32_to_str(0x231C4) // U+231C4 <cjk>
	0x5A: [`\u6659`].string() // U+6659 <cjk>
	0x5B: [`\u665A`].string() // U+665A <cjk>
	0x5C: [`\u6661`].string() // U+6661 <cjk>
	0x5D: [`\u6665`].string() // U+6665 <cjk>
	0x5E: [`\u6673`].string() // U+6673 <cjk>
	0x5F: [`\u6677`].string() // U+6677 <cjk>
	0x60: [`\u6678`].string() // U+6678 <cjk>
	0x61: [`\u668D`].string() // U+668D <cjk>
	0x62: [`\uFA43`].string() // U+FA43 CJK COMPATIBILITY IDEOGRAPH-FA43
	0x63: [`\u66A0`].string() // U+66A0 <cjk>
	0x64: [`\u66B2`].string() // U+66B2 <cjk>
	0x65: [`\u66BB`].string() // U+66BB <cjk>
	0x66: [`\u66C6`].string() // U+66C6 <cjk>
	0x67: [`\u66C8`].string() // U+66C8 <cjk>
	0x68: [`\u3B22`].string() // U+3B22 <cjk>
	0x69: [`\u66DB`].string() // U+66DB <cjk>
	0x6A: [`\u66E8`].string() // U+66E8 <cjk>
	0x6B: [`\u66FA`].string() // U+66FA <cjk>
	0x6C: [`\u6713`].string() // U+6713 <cjk>
	0x6D: [`\uF929`].string() // U+F929 CJK COMPATIBILITY IDEOGRAPH-F929
	0x6E: [`\u6733`].string() // U+6733 <cjk>
	0x6F: [`\u6766`].string() // U+6766 <cjk>
	0x70: [`\u6747`].string() // U+6747 <cjk>
	0x71: [`\u6748`].string() // U+6748 <cjk>
	0x72: [`\u677B`].string() // U+677B <cjk>
	0x73: [`\u6781`].string() // U+6781 <cjk>
	0x74: [`\u6793`].string() // U+6793 <cjk>
	0x75: [`\u6798`].string() // U+6798 <cjk>
	0x76: [`\u679B`].string() // U+679B <cjk>
	0x77: [`\u67BB`].string() // U+67BB <cjk>
	0x78: [`\u67F9`].string() // U+67F9 <cjk>
	0x79: [`\u67C0`].string() // U+67C0 <cjk>
	0x7A: [`\u67D7`].string() // U+67D7 <cjk>
	0x7B: [`\u67FC`].string() // U+67FC <cjk>
	0x7C: [`\u6801`].string() // U+6801 <cjk>
	0x7D: [`\u6852`].string() // U+6852 <cjk>
	0x7E: [`\u681D`].string() // U+681D <cjk>
	0x80: [`\u682C`].string() // U+682C <cjk>
	0x81: [`\u6831`].string() // U+6831 <cjk>
	0x82: [`\u685B`].string() // U+685B <cjk>
	0x83: [`\u6872`].string() // U+6872 <cjk>
	0x84: [`\u6875`].string() // U+6875 <cjk>
	0x85: [`\uFA44`].string() // U+FA44 CJK COMPATIBILITY IDEOGRAPH-FA44
	0x86: [`\u68A3`].string() // U+68A3 <cjk>
	0x87: [`\u68A5`].string() // U+68A5 <cjk>
	0x88: [`\u68B2`].string() // U+68B2 <cjk>
	0x89: [`\u68C8`].string() // U+68C8 <cjk>
	0x8A: [`\u68D0`].string() // U+68D0 <cjk>
	0x8B: [`\u68E8`].string() // U+68E8 <cjk>
	0x8C: [`\u68ED`].string() // U+68ED <cjk>
	0x8D: [`\u68F0`].string() // U+68F0 <cjk>
	0x8E: [`\u68F1`].string() // U+68F1 <cjk>
	0x8F: [`\u68FC`].string() // U+68FC <cjk>
	0x90: [`\u690A`].string() // U+690A <cjk>
	0x91: [`\u6949`].string() // U+6949 <cjk>
	0x92: utf32_to_str(0x235C4) // U+235C4 <cjk>
	0x93: [`\u6935`].string() // U+6935 <cjk>
	0x94: [`\u6942`].string() // U+6942 <cjk>
	0x95: [`\u6957`].string() // U+6957 <cjk>
	0x96: [`\u6963`].string() // U+6963 <cjk>
	0x97: [`\u6964`].string() // U+6964 <cjk>
	0x98: [`\u6968`].string() // U+6968 <cjk>
	0x99: [`\u6980`].string() // U+6980 <cjk>
	0x9A: [`\uFA14`].string() // U+FA14 CJK COMPATIBILITY IDEOGRAPH-FA14
	0x9B: [`\u69A5`].string() // U+69A5 <cjk>
	0x9C: [`\u69AD`].string() // U+69AD <cjk>
	0x9D: [`\u69CF`].string() // U+69CF <cjk>
	0x9E: [`\u3BB6`].string() // U+3BB6 <cjk>
	0x9F: [`\u3BC3`].string() // U+3BC3 <cjk>
	0xA0: [`\u69E2`].string() // U+69E2 <cjk>
	0xA1: [`\u69E9`].string() // U+69E9 <cjk>
	0xA2: [`\u69EA`].string() // U+69EA <cjk>
	0xA3: [`\u69F5`].string() // U+69F5 <cjk>
	0xA4: [`\u69F6`].string() // U+69F6 <cjk>
	0xA5: [`\u6A0F`].string() // U+6A0F <cjk>
	0xA6: [`\u6A15`].string() // U+6A15 <cjk>
	0xA7: utf32_to_str(0x2373F) // U+2373F <cjk>
	0xA8: [`\u6A3B`].string() // U+6A3B <cjk>
	0xA9: [`\u6A3E`].string() // U+6A3E <cjk>
	0xAA: [`\u6A45`].string() // U+6A45 <cjk>
	0xAB: [`\u6A50`].string() // U+6A50 <cjk>
	0xAC: [`\u6A56`].string() // U+6A56 <cjk>
	0xAD: [`\u6A5B`].string() // U+6A5B <cjk>
	0xAE: [`\u6A6B`].string() // U+6A6B <cjk>
	0xAF: [`\u6A73`].string() // U+6A73 <cjk>
	0xB0: utf32_to_str(0x23763) // U+23763 <cjk>
	0xB1: [`\u6A89`].string() // U+6A89 <cjk>
	0xB2: [`\u6A94`].string() // U+6A94 <cjk>
	0xB3: [`\u6A9D`].string() // U+6A9D <cjk>
	0xB4: [`\u6A9E`].string() // U+6A9E <cjk>
	0xB5: [`\u6AA5`].string() // U+6AA5 <cjk>
	0xB6: [`\u6AE4`].string() // U+6AE4 <cjk>
	0xB7: [`\u6AE7`].string() // U+6AE7 <cjk>
	0xB8: [`\u3C0F`].string() // U+3C0F <cjk>
	0xB9: [`\uF91D`].string() // U+F91D CJK COMPATIBILITY IDEOGRAPH-F91D
	0xBA: [`\u6B1B`].string() // U+6B1B <cjk>
	0xBB: [`\u6B1E`].string() // U+6B1E <cjk>
	0xBC: [`\u6B2C`].string() // U+6B2C <cjk>
	0xBD: [`\u6B35`].string() // U+6B35 <cjk>
	0xBE: [`\u6B46`].string() // U+6B46 <cjk>
	0xBF: [`\u6B56`].string() // U+6B56 <cjk>
	0xC0: [`\u6B60`].string() // U+6B60 <cjk>
	0xC1: [`\u6B65`].string() // U+6B65 <cjk>
	0xC2: [`\u6B67`].string() // U+6B67 <cjk>
	0xC3: [`\u6B77`].string() // U+6B77 <cjk>
	0xC4: [`\u6B82`].string() // U+6B82 <cjk>
	0xC5: [`\u6BA9`].string() // U+6BA9 <cjk>
	0xC6: [`\u6BAD`].string() // U+6BAD <cjk>
	0xC7: [`\uF970`].string() // U+F970 CJK COMPATIBILITY IDEOGRAPH-F970
	0xC8: [`\u6BCF`].string() // U+6BCF <cjk>
	0xC9: [`\u6BD6`].string() // U+6BD6 <cjk>
	0xCA: [`\u6BD7`].string() // U+6BD7 <cjk>
	0xCB: [`\u6BFF`].string() // U+6BFF <cjk>
	0xCC: [`\u6C05`].string() // U+6C05 <cjk>
	0xCD: [`\u6C10`].string() // U+6C10 <cjk>
	0xCE: [`\u6C33`].string() // U+6C33 <cjk>
	0xCF: [`\u6C59`].string() // U+6C59 <cjk>
	0xD0: [`\u6C5C`].string() // U+6C5C <cjk>
	0xD1: [`\u6CAA`].string() // U+6CAA <cjk>
	0xD2: [`\u6C74`].string() // U+6C74 <cjk>
	0xD3: [`\u6C76`].string() // U+6C76 <cjk>
	0xD4: [`\u6C85`].string() // U+6C85 <cjk>
	0xD5: [`\u6C86`].string() // U+6C86 <cjk>
	0xD6: [`\u6C98`].string() // U+6C98 <cjk>
	0xD7: [`\u6C9C`].string() // U+6C9C <cjk>
	0xD8: [`\u6CFB`].string() // U+6CFB <cjk>
	0xD9: [`\u6CC6`].string() // U+6CC6 <cjk>
	0xDA: [`\u6CD4`].string() // U+6CD4 <cjk>
	0xDB: [`\u6CE0`].string() // U+6CE0 <cjk>
	0xDC: [`\u6CEB`].string() // U+6CEB <cjk>
	0xDD: [`\u6CEE`].string() // U+6CEE <cjk>
	0xDE: utf32_to_str(0x23CFE) // U+23CFE <cjk>
	0xDF: [`\u6D04`].string() // U+6D04 <cjk>
	0xE0: [`\u6D0E`].string() // U+6D0E <cjk>
	0xE1: [`\u6D2E`].string() // U+6D2E <cjk>
	0xE2: [`\u6D31`].string() // U+6D31 <cjk>
	0xE3: [`\u6D39`].string() // U+6D39 <cjk>
	0xE4: [`\u6D3F`].string() // U+6D3F <cjk>
	0xE5: [`\u6D58`].string() // U+6D58 <cjk>
	0xE6: [`\u6D65`].string() // U+6D65 <cjk>
	0xE7: [`\uFA45`].string() // U+FA45 CJK COMPATIBILITY IDEOGRAPH-FA45
	0xE8: [`\u6D82`].string() // U+6D82 <cjk>
	0xE9: [`\u6D87`].string() // U+6D87 <cjk>
	0xEA: [`\u6D89`].string() // U+6D89 <cjk>
	0xEB: [`\u6D94`].string() // U+6D94 <cjk>
	0xEC: [`\u6DAA`].string() // U+6DAA <cjk>
	0xED: [`\u6DAC`].string() // U+6DAC <cjk>
	0xEE: [`\u6DBF`].string() // U+6DBF <cjk>
	0xEF: [`\u6DC4`].string() // U+6DC4 <cjk>
	0xF0: [`\u6DD6`].string() // U+6DD6 <cjk>
	0xF1: [`\u6DDA`].string() // U+6DDA <cjk>
	0xF2: [`\u6DDB`].string() // U+6DDB <cjk>
	0xF3: [`\u6DDD`].string() // U+6DDD <cjk>
	0xF4: [`\u6DFC`].string() // U+6DFC <cjk>
	0xF5: [`\uFA46`].string() // U+FA46 CJK COMPATIBILITY IDEOGRAPH-FA46
	0xF6: [`\u6E34`].string() // U+6E34 <cjk>
	0xF7: [`\u6E44`].string() // U+6E44 <cjk>
	0xF8: [`\u6E5C`].string() // U+6E5C <cjk>
	0xF9: [`\u6E5E`].string() // U+6E5E <cjk>
	0xFA: [`\u6EAB`].string() // U+6EAB <cjk>
	0xFB: [`\u6EB1`].string() // U+6EB1 <cjk>
	0xFC: [`\u6EC1`].string() // U+6EC1 <cjk>
}

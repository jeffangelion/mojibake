module mojibake

const jis_x_0213_doublebyte_0x9e = {
	0x40: [`\u66C4`].string() // U+66C4 <cjk>
	0x41: [`\u66B8`].string() // U+66B8 <cjk>
	0x42: [`\u66D6`].string() // U+66D6 <cjk>
	0x43: [`\u66DA`].string() // U+66DA <cjk>
	0x44: [`\u66E0`].string() // U+66E0 <cjk>
	0x45: [`\u663F`].string() // U+663F <cjk>
	0x46: [`\u66E6`].string() // U+66E6 <cjk>
	0x47: [`\u66E9`].string() // U+66E9 <cjk>
	0x48: [`\u66F0`].string() // U+66F0 <cjk>
	0x49: [`\u66F5`].string() // U+66F5 <cjk>
	0x4A: [`\u66F7`].string() // U+66F7 <cjk>
	0x4B: [`\u670F`].string() // U+670F <cjk>
	0x4C: [`\u6716`].string() // U+6716 <cjk>
	0x4D: [`\u671E`].string() // U+671E <cjk>
	0x4E: [`\u6726`].string() // U+6726 <cjk>
	0x4F: [`\u6727`].string() // U+6727 <cjk>
	0x50: [`\u9738`].string() // U+9738 <cjk>
	0x51: [`\u672E`].string() // U+672E <cjk>
	0x52: [`\u673F`].string() // U+673F <cjk>
	0x53: [`\u6736`].string() // U+6736 <cjk>
	0x54: [`\u6741`].string() // U+6741 <cjk>
	0x55: [`\u6738`].string() // U+6738 <cjk>
	0x56: [`\u6737`].string() // U+6737 <cjk>
	0x57: [`\u6746`].string() // U+6746 <cjk>
	0x58: [`\u675E`].string() // U+675E <cjk>
	0x59: [`\u6760`].string() // U+6760 <cjk>
	0x5A: [`\u6759`].string() // U+6759 <cjk>
	0x5B: [`\u6763`].string() // U+6763 <cjk>
	0x5C: [`\u6764`].string() // U+6764 <cjk>
	0x5D: [`\u6789`].string() // U+6789 <cjk>
	0x5E: [`\u6770`].string() // U+6770 <cjk>
	0x5F: [`\u67A9`].string() // U+67A9 <cjk>
	0x60: [`\u677C`].string() // U+677C <cjk>
	0x61: [`\u676A`].string() // U+676A <cjk>
	0x62: [`\u678C`].string() // U+678C <cjk>
	0x63: [`\u678B`].string() // U+678B <cjk>
	0x64: [`\u67A6`].string() // U+67A6 <cjk>
	0x65: [`\u67A1`].string() // U+67A1 <cjk>
	0x66: [`\u6785`].string() // U+6785 <cjk>
	0x67: [`\u67B7`].string() // U+67B7 <cjk>
	0x68: [`\u67EF`].string() // U+67EF <cjk>
	0x69: [`\u67B4`].string() // U+67B4 <cjk>
	0x6A: [`\u67EC`].string() // U+67EC <cjk>
	0x6B: [`\u67B3`].string() // U+67B3 <cjk>
	0x6C: [`\u67E9`].string() // U+67E9 <cjk>
	0x6D: [`\u67B8`].string() // U+67B8 <cjk>
	0x6E: [`\u67E4`].string() // U+67E4 <cjk>
	0x6F: [`\u67DE`].string() // U+67DE <cjk>
	0x70: [`\u67DD`].string() // U+67DD <cjk>
	0x71: [`\u67E2`].string() // U+67E2 <cjk>
	0x72: [`\u67EE`].string() // U+67EE <cjk>
	0x73: [`\u67B9`].string() // U+67B9 <cjk>
	0x74: [`\u67CE`].string() // U+67CE <cjk>
	0x75: [`\u67C6`].string() // U+67C6 <cjk>
	0x76: [`\u67E7`].string() // U+67E7 <cjk>
	0x77: [`\u6A9C`].string() // U+6A9C <cjk>
	0x78: [`\u681E`].string() // U+681E <cjk>
	0x79: [`\u6846`].string() // U+6846 <cjk>
	0x7A: [`\u6829`].string() // U+6829 <cjk>
	0x7B: [`\u6840`].string() // U+6840 <cjk>
	0x7C: [`\u684D`].string() // U+684D <cjk>
	0x7D: [`\u6832`].string() // U+6832 <cjk>
	0x7E: [`\u684E`].string() // U+684E <cjk>
	0x80: [`\u68B3`].string() // U+68B3 <cjk>
	0x81: [`\u682B`].string() // U+682B <cjk>
	0x82: [`\u6859`].string() // U+6859 <cjk>
	0x83: [`\u6863`].string() // U+6863 <cjk>
	0x84: [`\u6877`].string() // U+6877 <cjk>
	0x85: [`\u687F`].string() // U+687F <cjk>
	0x86: [`\u689F`].string() // U+689F <cjk>
	0x87: [`\u688F`].string() // U+688F <cjk>
	0x88: [`\u68AD`].string() // U+68AD <cjk>
	0x89: [`\u6894`].string() // U+6894 <cjk>
	0x8A: [`\u689D`].string() // U+689D <cjk>
	0x8B: [`\u689B`].string() // U+689B <cjk>
	0x8C: [`\u6883`].string() // U+6883 <cjk>
	0x8D: [`\u6AAE`].string() // U+6AAE <cjk>
	0x8E: [`\u68B9`].string() // U+68B9 <cjk>
	0x8F: [`\u6874`].string() // U+6874 <cjk>
	0x90: [`\u68B5`].string() // U+68B5 <cjk>
	0x91: [`\u68A0`].string() // U+68A0 <cjk>
	0x92: [`\u68BA`].string() // U+68BA <cjk>
	0x93: [`\u690F`].string() // U+690F <cjk>
	0x94: [`\u688D`].string() // U+688D <cjk>
	0x95: [`\u687E`].string() // U+687E <cjk>
	0x96: [`\u6901`].string() // U+6901 <cjk>
	0x97: [`\u68CA`].string() // U+68CA <cjk>
	0x98: [`\u6908`].string() // U+6908 <cjk>
	0x99: [`\u68D8`].string() // U+68D8 <cjk>
	0x9A: [`\u6922`].string() // U+6922 <cjk>
	0x9B: [`\u6926`].string() // U+6926 <cjk>
	0x9C: [`\u68E1`].string() // U+68E1 <cjk>
	0x9D: [`\u690C`].string() // U+690C <cjk>
	0x9E: [`\u68CD`].string() // U+68CD <cjk>
	0x9F: [`\u68D4`].string() // U+68D4 <cjk>
	0xA0: [`\u68E7`].string() // U+68E7 <cjk>
	0xA1: [`\u68D5`].string() // U+68D5 <cjk>
	0xA2: [`\u6936`].string() // U+6936 <cjk>
	0xA3: [`\u6912`].string() // U+6912 <cjk>
	0xA4: [`\u6904`].string() // U+6904 <cjk>
	0xA5: [`\u68D7`].string() // U+68D7 <cjk>
	0xA6: [`\u68E3`].string() // U+68E3 <cjk>
	0xA7: [`\u6925`].string() // U+6925 <cjk>
	0xA8: [`\u68F9`].string() // U+68F9 <cjk>
	0xA9: [`\u68E0`].string() // U+68E0 <cjk>
	0xAA: [`\u68EF`].string() // U+68EF <cjk>
	0xAB: [`\u6928`].string() // U+6928 <cjk>
	0xAC: [`\u692A`].string() // U+692A <cjk>
	0xAD: [`\u691A`].string() // U+691A <cjk>
	0xAE: [`\u6923`].string() // U+6923 <cjk>
	0xAF: [`\u6921`].string() // U+6921 <cjk>
	0xB0: [`\u68C6`].string() // U+68C6 <cjk>
	0xB1: [`\u6979`].string() // U+6979 <cjk>
	0xB2: [`\u6977`].string() // U+6977 <cjk>
	0xB3: [`\u695C`].string() // U+695C <cjk>
	0xB4: [`\u6978`].string() // U+6978 <cjk>
	0xB5: [`\u696B`].string() // U+696B <cjk>
	0xB6: [`\u6954`].string() // U+6954 <cjk>
	0xB7: [`\u697E`].string() // U+697E <cjk>
	0xB8: [`\u696E`].string() // U+696E <cjk>
	0xB9: [`\u6939`].string() // U+6939 <cjk>
	0xBA: [`\u6974`].string() // U+6974 <cjk>
	0xBB: [`\u693D`].string() // U+693D <cjk>
	0xBC: [`\u6959`].string() // U+6959 <cjk>
	0xBD: [`\u6930`].string() // U+6930 <cjk>
	0xBE: [`\u6961`].string() // U+6961 <cjk>
	0xBF: [`\u695E`].string() // U+695E <cjk>
	0xC0: [`\u695D`].string() // U+695D <cjk>
	0xC1: [`\u6981`].string() // U+6981 <cjk>
	0xC2: [`\u696A`].string() // U+696A <cjk>
	0xC3: [`\u69B2`].string() // U+69B2 <cjk>
	0xC4: [`\u69AE`].string() // U+69AE <cjk>
	0xC5: [`\u69D0`].string() // U+69D0 <cjk>
	0xC6: [`\u69BF`].string() // U+69BF <cjk>
	0xC7: [`\u69C1`].string() // U+69C1 <cjk>
	0xC8: [`\u69D3`].string() // U+69D3 <cjk>
	0xC9: [`\u69BE`].string() // U+69BE <cjk>
	0xCA: [`\u69CE`].string() // U+69CE <cjk>
	0xCB: [`\u5BE8`].string() // U+5BE8 <cjk>
	0xCC: [`\u69CA`].string() // U+69CA <cjk>
	0xCD: [`\u69DD`].string() // U+69DD <cjk>
	0xCE: [`\u69BB`].string() // U+69BB <cjk>
	0xCF: [`\u69C3`].string() // U+69C3 <cjk>
	0xD0: [`\u69A7`].string() // U+69A7 <cjk>
	0xD1: [`\u6A2E`].string() // U+6A2E <cjk>
	0xD2: [`\u6991`].string() // U+6991 <cjk>
	0xD3: [`\u69A0`].string() // U+69A0 <cjk>
	0xD4: [`\u699C`].string() // U+699C <cjk>
	0xD5: [`\u6995`].string() // U+6995 <cjk>
	0xD6: [`\u69B4`].string() // U+69B4 <cjk>
	0xD7: [`\u69DE`].string() // U+69DE <cjk>
	0xD8: [`\u69E8`].string() // U+69E8 <cjk>
	0xD9: [`\u6A02`].string() // U+6A02 <cjk>
	0xDA: [`\u6A1B`].string() // U+6A1B <cjk>
	0xDB: [`\u69FF`].string() // U+69FF <cjk>
	0xDC: [`\u6B0A`].string() // U+6B0A <cjk>
	0xDD: [`\u69F9`].string() // U+69F9 <cjk>
	0xDE: [`\u69F2`].string() // U+69F2 <cjk>
	0xDF: [`\u69E7`].string() // U+69E7 <cjk>
	0xE0: [`\u6A05`].string() // U+6A05 <cjk>
	0xE1: [`\u69B1`].string() // U+69B1 <cjk>
	0xE2: [`\u6A1E`].string() // U+6A1E <cjk>
	0xE3: [`\u69ED`].string() // U+69ED <cjk>
	0xE4: [`\u6A14`].string() // U+6A14 <cjk>
	0xE5: [`\u69EB`].string() // U+69EB <cjk>
	0xE6: [`\u6A0A`].string() // U+6A0A <cjk>
	0xE7: [`\u6A12`].string() // U+6A12 <cjk>
	0xE8: [`\u6AC1`].string() // U+6AC1 <cjk>
	0xE9: [`\u6A23`].string() // U+6A23 <cjk>
	0xEA: [`\u6A13`].string() // U+6A13 <cjk>
	0xEB: [`\u6A44`].string() // U+6A44 <cjk>
	0xEC: [`\u6A0C`].string() // U+6A0C <cjk>
	0xED: [`\u6A72`].string() // U+6A72 <cjk>
	0xEE: [`\u6A36`].string() // U+6A36 <cjk>
	0xEF: [`\u6A78`].string() // U+6A78 <cjk>
	0xF0: [`\u6A47`].string() // U+6A47 <cjk>
	0xF1: [`\u6A62`].string() // U+6A62 <cjk>
	0xF2: [`\u6A59`].string() // U+6A59 <cjk>
	0xF3: [`\u6A66`].string() // U+6A66 <cjk>
	0xF4: [`\u6A48`].string() // U+6A48 <cjk>
	0xF5: [`\u6A38`].string() // U+6A38 <cjk>
	0xF6: [`\u6A22`].string() // U+6A22 <cjk>
	0xF7: [`\u6A90`].string() // U+6A90 <cjk>
	0xF8: [`\u6A8D`].string() // U+6A8D <cjk>
	0xF9: [`\u6AA0`].string() // U+6AA0 <cjk>
	0xFA: [`\u6A84`].string() // U+6A84 <cjk>
	0xFB: [`\u6AA2`].string() // U+6AA2 <cjk>
	0xFC: [`\u6AA3`].string() // U+6AA3 <cjk>
}

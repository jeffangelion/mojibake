module mojibake

const jis_x_0213_doublebyte_0xfb = {
	0x40: utf32_to_str(0x28A29) // U+28A29 <cjk>
	0x41: [`\u92F7`].string() // U+92F7 <cjk>
	0x42: [`\u92F9`].string() // U+92F9 <cjk>
	0x43: [`\u92FB`].string() // U+92FB <cjk>
	0x44: [`\u9302`].string() // U+9302 <cjk>
	0x45: [`\u930D`].string() // U+930D <cjk>
	0x46: [`\u9315`].string() // U+9315 <cjk>
	0x47: [`\u931D`].string() // U+931D <cjk>
	0x48: [`\u931E`].string() // U+931E <cjk>
	0x49: [`\u9327`].string() // U+9327 <cjk>
	0x4A: [`\u9329`].string() // U+9329 <cjk>
	0x4B: utf32_to_str(0x28A71) // U+28A71 <cjk>
	0x4C: utf32_to_str(0x28A43) // U+28A43 <cjk>
	0x4D: [`\u9347`].string() // U+9347 <cjk>
	0x4E: [`\u9351`].string() // U+9351 <cjk>
	0x4F: [`\u9357`].string() // U+9357 <cjk>
	0x50: [`\u935A`].string() // U+935A <cjk>
	0x51: [`\u936B`].string() // U+936B <cjk>
	0x52: [`\u9371`].string() // U+9371 <cjk>
	0x53: [`\u9373`].string() // U+9373 <cjk>
	0x54: [`\u93A1`].string() // U+93A1 <cjk>
	0x55: utf32_to_str(0x28A99) // U+28A99 <cjk>
	0x56: utf32_to_str(0x28ACD) // U+28ACD <cjk>
	0x57: [`\u9388`].string() // U+9388 <cjk>
	0x58: [`\u938B`].string() // U+938B <cjk>
	0x59: [`\u938F`].string() // U+938F <cjk>
	0x5A: [`\u939E`].string() // U+939E <cjk>
	0x5B: [`\u93F5`].string() // U+93F5 <cjk>
	0x5C: utf32_to_str(0x28AE4) // U+28AE4 <cjk>
	0x5D: utf32_to_str(0x28ADD) // U+28ADD <cjk>
	0x5E: [`\u93F1`].string() // U+93F1 <cjk>
	0x5F: [`\u93C1`].string() // U+93C1 <cjk>
	0x60: [`\u93C7`].string() // U+93C7 <cjk>
	0x61: [`\u93DC`].string() // U+93DC <cjk>
	0x62: [`\u93E2`].string() // U+93E2 <cjk>
	0x63: [`\u93E7`].string() // U+93E7 <cjk>
	0x64: [`\u9409`].string() // U+9409 <cjk>
	0x65: [`\u940F`].string() // U+940F <cjk>
	0x66: [`\u9416`].string() // U+9416 <cjk>
	0x67: [`\u9417`].string() // U+9417 <cjk>
	0x68: [`\u93FB`].string() // U+93FB <cjk>
	0x69: [`\u9432`].string() // U+9432 <cjk>
	0x6A: [`\u9434`].string() // U+9434 <cjk>
	0x6B: [`\u943B`].string() // U+943B <cjk>
	0x6C: [`\u9445`].string() // U+9445 <cjk>
	0x6D: utf32_to_str(0x28BC1) // U+28BC1 <cjk>
	0x6E: utf32_to_str(0x28BEF) // U+28BEF <cjk>
	0x6F: [`\u946D`].string() // U+946D <cjk>
	0x70: [`\u946F`].string() // U+946F <cjk>
	0x71: [`\u9578`].string() // U+9578 <cjk>
	0x72: [`\u9579`].string() // U+9579 <cjk>
	0x73: [`\u9586`].string() // U+9586 <cjk>
	0x74: [`\u958C`].string() // U+958C <cjk>
	0x75: [`\u958D`].string() // U+958D <cjk>
	0x76: utf32_to_str(0x28D10) // U+28D10 <cjk>
	0x77: [`\u95AB`].string() // U+95AB <cjk>
	0x78: [`\u95B4`].string() // U+95B4 <cjk>
	0x79: utf32_to_str(0x28D71) // U+28D71 <cjk>
	0x7A: [`\u95C8`].string() // U+95C8 <cjk>
	0x7B: utf32_to_str(0x28DFB) // U+28DFB <cjk>
	0x7C: utf32_to_str(0x28E1F) // U+28E1F <cjk>
	0x7D: [`\u962C`].string() // U+962C <cjk>
	0x7E: [`\u9633`].string() // U+9633 <cjk>
	0x80: [`\u9634`].string() // U+9634 <cjk>
	0x81: utf32_to_str(0x28E36) // U+28E36 <cjk>
	0x82: [`\u963C`].string() // U+963C <cjk>
	0x83: [`\u9641`].string() // U+9641 <cjk>
	0x84: [`\u9661`].string() // U+9661 <cjk>
	0x85: utf32_to_str(0x28E89) // U+28E89 <cjk>
	0x86: [`\u9682`].string() // U+9682 <cjk>
	0x87: utf32_to_str(0x28EEB) // U+28EEB <cjk>
	0x88: [`\u969A`].string() // U+969A <cjk>
	0x89: utf32_to_str(0x28F32) // U+28F32 <cjk>
	0x8A: [`\u49E7`].string() // U+49E7 <cjk>
	0x8B: [`\u96A9`].string() // U+96A9 <cjk>
	0x8C: [`\u96AF`].string() // U+96AF <cjk>
	0x8D: [`\u96B3`].string() // U+96B3 <cjk>
	0x8E: [`\u96BA`].string() // U+96BA <cjk>
	0x8F: [`\u96BD`].string() // U+96BD <cjk>
	0x90: [`\u49FA`].string() // U+49FA <cjk>
	0x91: utf32_to_str(0x28FF8) // U+28FF8 <cjk>
	0x92: [`\u96D8`].string() // U+96D8 <cjk>
	0x93: [`\u96DA`].string() // U+96DA <cjk>
	0x94: [`\u96DD`].string() // U+96DD <cjk>
	0x95: [`\u4A04`].string() // U+4A04 <cjk>
	0x96: [`\u9714`].string() // U+9714 <cjk>
	0x97: [`\u9723`].string() // U+9723 <cjk>
	0x98: [`\u4A29`].string() // U+4A29 <cjk>
	0x99: [`\u9736`].string() // U+9736 <cjk>
	0x9A: [`\u9741`].string() // U+9741 <cjk>
	0x9B: [`\u9747`].string() // U+9747 <cjk>
	0x9C: [`\u9755`].string() // U+9755 <cjk>
	0x9D: [`\u9757`].string() // U+9757 <cjk>
	0x9E: [`\u975B`].string() // U+975B <cjk>
	0x9F: [`\u976A`].string() // U+976A <cjk>
	0xA0: utf32_to_str(0x292A0) // U+292A0 <cjk>
	0xA1: utf32_to_str(0x292B1) // U+292B1 <cjk>
	0xA2: [`\u9796`].string() // U+9796 <cjk>
	0xA3: [`\u979A`].string() // U+979A <cjk>
	0xA4: [`\u979E`].string() // U+979E <cjk>
	0xA5: [`\u97A2`].string() // U+97A2 <cjk>
	0xA6: [`\u97B1`].string() // U+97B1 <cjk>
	0xA7: [`\u97B2`].string() // U+97B2 <cjk>
	0xA8: [`\u97BE`].string() // U+97BE <cjk>
	0xA9: [`\u97CC`].string() // U+97CC <cjk>
	0xAA: [`\u97D1`].string() // U+97D1 <cjk>
	0xAB: [`\u97D4`].string() // U+97D4 <cjk>
	0xAC: [`\u97D8`].string() // U+97D8 <cjk>
	0xAD: [`\u97D9`].string() // U+97D9 <cjk>
	0xAE: [`\u97E1`].string() // U+97E1 <cjk>
	0xAF: [`\u97F1`].string() // U+97F1 <cjk>
	0xB0: [`\u9804`].string() // U+9804 <cjk>
	0xB1: [`\u980D`].string() // U+980D <cjk>
	0xB2: [`\u980E`].string() // U+980E <cjk>
	0xB3: [`\u9814`].string() // U+9814 <cjk>
	0xB4: [`\u9816`].string() // U+9816 <cjk>
	0xB5: [`\u4ABC`].string() // U+4ABC <cjk>
	0xB6: utf32_to_str(0x29490) // U+29490 <cjk>
	0xB7: [`\u9823`].string() // U+9823 <cjk>
	0xB8: [`\u9832`].string() // U+9832 <cjk>
	0xB9: [`\u9833`].string() // U+9833 <cjk>
	0xBA: [`\u9825`].string() // U+9825 <cjk>
	0xBB: [`\u9847`].string() // U+9847 <cjk>
	0xBC: [`\u9866`].string() // U+9866 <cjk>
	0xBD: [`\u98AB`].string() // U+98AB <cjk>
	0xBE: [`\u98AD`].string() // U+98AD <cjk>
	0xBF: [`\u98B0`].string() // U+98B0 <cjk>
	0xC0: utf32_to_str(0x295CF) // U+295CF <cjk>
	0xC1: [`\u98B7`].string() // U+98B7 <cjk>
	0xC2: [`\u98B8`].string() // U+98B8 <cjk>
	0xC3: [`\u98BB`].string() // U+98BB <cjk>
	0xC4: [`\u98BC`].string() // U+98BC <cjk>
	0xC5: [`\u98BF`].string() // U+98BF <cjk>
	0xC6: [`\u98C2`].string() // U+98C2 <cjk>
	0xC7: [`\u98C7`].string() // U+98C7 <cjk>
	0xC8: [`\u98CB`].string() // U+98CB <cjk>
	0xC9: [`\u98E0`].string() // U+98E0 <cjk>
	0xCA: utf32_to_str(0x2967F) // U+2967F <cjk>
	0xCB: [`\u98E1`].string() // U+98E1 <cjk>
	0xCC: [`\u98E3`].string() // U+98E3 <cjk>
	0xCD: [`\u98E5`].string() // U+98E5 <cjk>
	0xCE: [`\u98EA`].string() // U+98EA <cjk>
	0xCF: [`\u98F0`].string() // U+98F0 <cjk>
	0xD0: [`\u98F1`].string() // U+98F1 <cjk>
	0xD1: [`\u98F3`].string() // U+98F3 <cjk>
	0xD2: [`\u9908`].string() // U+9908 <cjk>
	0xD3: [`\u4B3B`].string() // U+4B3B <cjk>
	0xD4: utf32_to_str(0x296F0) // U+296F0 <cjk>
	0xD5: [`\u9916`].string() // U+9916 <cjk>
	0xD6: [`\u9917`].string() // U+9917 <cjk>
	0xD7: utf32_to_str(0x29719) // U+29719 <cjk>
	0xD8: [`\u991A`].string() // U+991A <cjk>
	0xD9: [`\u991B`].string() // U+991B <cjk>
	0xDA: [`\u991C`].string() // U+991C <cjk>
	0xDB: utf32_to_str(0x29750) // U+29750 <cjk>
	0xDC: [`\u9931`].string() // U+9931 <cjk>
	0xDD: [`\u9932`].string() // U+9932 <cjk>
	0xDE: [`\u9933`].string() // U+9933 <cjk>
	0xDF: [`\u993A`].string() // U+993A <cjk>
	0xE0: [`\u993B`].string() // U+993B <cjk>
	0xE1: [`\u993C`].string() // U+993C <cjk>
	0xE2: [`\u9940`].string() // U+9940 <cjk>
	0xE3: [`\u9941`].string() // U+9941 <cjk>
	0xE4: [`\u9946`].string() // U+9946 <cjk>
	0xE5: [`\u994D`].string() // U+994D <cjk>
	0xE6: [`\u994E`].string() // U+994E <cjk>
	0xE7: [`\u995C`].string() // U+995C <cjk>
	0xE8: [`\u995F`].string() // U+995F <cjk>
	0xE9: [`\u9960`].string() // U+9960 <cjk>
	0xEA: [`\u99A3`].string() // U+99A3 <cjk>
	0xEB: [`\u99A6`].string() // U+99A6 <cjk>
	0xEC: [`\u99B9`].string() // U+99B9 <cjk>
	0xED: [`\u99BD`].string() // U+99BD <cjk>
	0xEE: [`\u99BF`].string() // U+99BF <cjk>
	0xEF: [`\u99C3`].string() // U+99C3 <cjk>
	0xF0: [`\u99C9`].string() // U+99C9 <cjk>
	0xF1: [`\u99D4`].string() // U+99D4 <cjk>
	0xF2: [`\u99D9`].string() // U+99D9 <cjk>
	0xF3: [`\u99DE`].string() // U+99DE <cjk>
	0xF4: utf32_to_str(0x298C6) // U+298C6 <cjk>
	0xF5: [`\u99F0`].string() // U+99F0 <cjk>
	0xF6: [`\u99F9`].string() // U+99F9 <cjk>
	0xF7: [`\u99FC`].string() // U+99FC <cjk>
	0xF8: [`\u9A0A`].string() // U+9A0A <cjk>
	0xF9: [`\u9A11`].string() // U+9A11 <cjk>
	0xFA: [`\u9A16`].string() // U+9A16 <cjk>
	0xFB: [`\u9A1A`].string() // U+9A1A <cjk>
	0xFC: [`\u9A20`].string() // U+9A20 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x92 = {
	0x40: [`\u53E9`].string() // U+53E9 <cjk>
	0x41: [`\u4F46`].string() // U+4F46 <cjk>
	0x42: [`\u9054`].string() // U+9054 <cjk>
	0x43: [`\u8FB0`].string() // U+8FB0 <cjk>
	0x44: [`\u596A`].string() // U+596A <cjk>
	0x45: [`\u8131`].string() // U+8131 <cjk>
	0x46: [`\u5DFD`].string() // U+5DFD <cjk>
	0x47: [`\u7AEA`].string() // U+7AEA <cjk>
	0x48: [`\u8FBF`].string() // U+8FBF <cjk>
	0x49: [`\u68DA`].string() // U+68DA <cjk>
	0x4A: [`\u8C37`].string() // U+8C37 <cjk>
	0x4B: [`\u72F8`].string() // U+72F8 <cjk>
	0x4C: [`\u9C48`].string() // U+9C48 <cjk>
	0x4D: [`\u6A3D`].string() // U+6A3D <cjk>
	0x4E: [`\u8AB0`].string() // U+8AB0 <cjk>
	0x4F: [`\u4E39`].string() // U+4E39 <cjk>
	0x50: [`\u5358`].string() // U+5358 <cjk>
	0x51: [`\u5606`].string() // U+5606 <cjk>
	0x52: [`\u5766`].string() // U+5766 <cjk>
	0x53: [`\u62C5`].string() // U+62C5 <cjk>
	0x54: [`\u63A2`].string() // U+63A2 <cjk>
	0x55: [`\u65E6`].string() // U+65E6 <cjk>
	0x56: [`\u6B4E`].string() // U+6B4E <cjk>
	0x57: [`\u6DE1`].string() // U+6DE1 <cjk>
	0x58: [`\u6E5B`].string() // U+6E5B <cjk>
	0x59: [`\u70AD`].string() // U+70AD <cjk>
	0x5A: [`\u77ED`].string() // U+77ED <cjk>
	0x5B: [`\u7AEF`].string() // U+7AEF <cjk>
	0x5C: [`\u7BAA`].string() // U+7BAA <cjk>
	0x5D: [`\u7DBB`].string() // U+7DBB <cjk>
	0x5E: [`\u803D`].string() // U+803D <cjk>
	0x5F: [`\u80C6`].string() // U+80C6 <cjk>
	0x60: [`\u86CB`].string() // U+86CB <cjk>
	0x61: [`\u8A95`].string() // U+8A95 <cjk>
	0x62: [`\u935B`].string() // U+935B <cjk>
	0x63: [`\u56E3`].string() // U+56E3 <cjk>
	0x64: [`\u58C7`].string() // U+58C7 <cjk>
	0x65: [`\u5F3E`].string() // U+5F3E <cjk>
	0x66: [`\u65AD`].string() // U+65AD <cjk>
	0x67: [`\u6696`].string() // U+6696 <cjk>
	0x68: [`\u6A80`].string() // U+6A80 <cjk>
	0x69: [`\u6BB5`].string() // U+6BB5 <cjk>
	0x6A: [`\u7537`].string() // U+7537 <cjk>
	0x6B: [`\u8AC7`].string() // U+8AC7 <cjk>
	0x6C: [`\u5024`].string() // U+5024 <cjk>
	0x6D: [`\u77E5`].string() // U+77E5 <cjk>
	0x6E: [`\u5730`].string() // U+5730 <cjk>
	0x6F: [`\u5F1B`].string() // U+5F1B <cjk>
	0x70: [`\u6065`].string() // U+6065 <cjk>
	0x71: [`\u667A`].string() // U+667A <cjk>
	0x72: [`\u6C60`].string() // U+6C60 <cjk>
	0x73: [`\u75F4`].string() // U+75F4 <cjk>
	0x74: [`\u7A1A`].string() // U+7A1A <cjk>
	0x75: [`\u7F6E`].string() // U+7F6E <cjk>
	0x76: [`\u81F4`].string() // U+81F4 <cjk>
	0x77: [`\u8718`].string() // U+8718 <cjk>
	0x78: [`\u9045`].string() // U+9045 <cjk>
	0x79: [`\u99B3`].string() // U+99B3 <cjk>
	0x7A: [`\u7BC9`].string() // U+7BC9 <cjk>
	0x7B: [`\u755C`].string() // U+755C <cjk>
	0x7C: [`\u7AF9`].string() // U+7AF9 <cjk>
	0x7D: [`\u7B51`].string() // U+7B51 <cjk>
	0x7E: [`\u84C4`].string() // U+84C4 <cjk>
	0x80: [`\u9010`].string() // U+9010 <cjk>
	0x81: [`\u79E9`].string() // U+79E9 <cjk>
	0x82: [`\u7A92`].string() // U+7A92 <cjk>
	0x83: [`\u8336`].string() // U+8336 <cjk>
	0x84: [`\u5AE1`].string() // U+5AE1 <cjk>
	0x85: [`\u7740`].string() // U+7740 <cjk>
	0x86: [`\u4E2D`].string() // U+4E2D <cjk>
	0x87: [`\u4EF2`].string() // U+4EF2 <cjk>
	0x88: [`\u5B99`].string() // U+5B99 <cjk>
	0x89: [`\u5FE0`].string() // U+5FE0 <cjk>
	0x8A: [`\u62BD`].string() // U+62BD <cjk>
	0x8B: [`\u663C`].string() // U+663C <cjk>
	0x8C: [`\u67F1`].string() // U+67F1 <cjk>
	0x8D: [`\u6CE8`].string() // U+6CE8 <cjk>
	0x8E: [`\u866B`].string() // U+866B <cjk>
	0x8F: [`\u8877`].string() // U+8877 <cjk>
	0x90: [`\u8A3B`].string() // U+8A3B <cjk>
	0x91: [`\u914E`].string() // U+914E <cjk>
	0x92: [`\u92F3`].string() // U+92F3 <cjk>
	0x93: [`\u99D0`].string() // U+99D0 <cjk>
	0x94: [`\u6A17`].string() // U+6A17 <cjk>
	0x95: [`\u7026`].string() // U+7026 <cjk>
	0x96: [`\u732A`].string() // U+732A <cjk>
	0x97: [`\u82E7`].string() // U+82E7 <cjk>
	0x98: [`\u8457`].string() // U+8457 <cjk>
	0x99: [`\u8CAF`].string() // U+8CAF <cjk>
	0x9A: [`\u4E01`].string() // U+4E01 <cjk>
	0x9B: [`\u5146`].string() // U+5146 <cjk>
	0x9C: [`\u51CB`].string() // U+51CB <cjk>
	0x9D: [`\u558B`].string() // U+558B <cjk>
	0x9E: [`\u5BF5`].string() // U+5BF5 <cjk>
	0x9F: [`\u5E16`].string() // U+5E16 <cjk>
	0xA0: [`\u5E33`].string() // U+5E33 <cjk>
	0xA1: [`\u5E81`].string() // U+5E81 <cjk>
	0xA2: [`\u5F14`].string() // U+5F14 <cjk>
	0xA3: [`\u5F35`].string() // U+5F35 <cjk>
	0xA4: [`\u5F6B`].string() // U+5F6B <cjk>
	0xA5: [`\u5FB4`].string() // U+5FB4 <cjk>
	0xA6: [`\u61F2`].string() // U+61F2 <cjk>
	0xA7: [`\u6311`].string() // U+6311 <cjk>
	0xA8: [`\u66A2`].string() // U+66A2 <cjk>
	0xA9: [`\u671D`].string() // U+671D <cjk>
	0xAA: [`\u6F6E`].string() // U+6F6E <cjk>
	0xAB: [`\u7252`].string() // U+7252 <cjk>
	0xAC: [`\u753A`].string() // U+753A <cjk>
	0xAD: [`\u773A`].string() // U+773A <cjk>
	0xAE: [`\u8074`].string() // U+8074 <cjk>
	0xAF: [`\u8139`].string() // U+8139 <cjk>
	0xB0: [`\u8178`].string() // U+8178 <cjk>
	0xB1: [`\u8776`].string() // U+8776 <cjk>
	0xB2: [`\u8ABF`].string() // U+8ABF <cjk>
	0xB3: [`\u8ADC`].string() // U+8ADC <cjk>
	0xB4: [`\u8D85`].string() // U+8D85 <cjk>
	0xB5: [`\u8DF3`].string() // U+8DF3 <cjk>
	0xB6: [`\u929A`].string() // U+929A <cjk>
	0xB7: [`\u9577`].string() // U+9577 <cjk>
	0xB8: [`\u9802`].string() // U+9802 <cjk>
	0xB9: [`\u9CE5`].string() // U+9CE5 <cjk>
	0xBA: [`\u52C5`].string() // U+52C5 <cjk>
	0xBB: [`\u6357`].string() // U+6357 <cjk>
	0xBC: [`\u76F4`].string() // U+76F4 <cjk>
	0xBD: [`\u6715`].string() // U+6715 <cjk>
	0xBE: [`\u6C88`].string() // U+6C88 <cjk>
	0xBF: [`\u73CD`].string() // U+73CD <cjk>
	0xC0: [`\u8CC3`].string() // U+8CC3 <cjk>
	0xC1: [`\u93AE`].string() // U+93AE <cjk>
	0xC2: [`\u9673`].string() // U+9673 <cjk>
	0xC3: [`\u6D25`].string() // U+6D25 <cjk>
	0xC4: [`\u589C`].string() // U+589C <cjk>
	0xC5: [`\u690E`].string() // U+690E <cjk>
	0xC6: [`\u69CC`].string() // U+69CC <cjk>
	0xC7: [`\u8FFD`].string() // U+8FFD <cjk>
	0xC8: [`\u939A`].string() // U+939A <cjk>
	0xC9: [`\u75DB`].string() // U+75DB <cjk>
	0xCA: [`\u901A`].string() // U+901A <cjk>
	0xCB: [`\u585A`].string() // U+585A <cjk>
	0xCC: [`\u6802`].string() // U+6802 <cjk>
	0xCD: [`\u63B4`].string() // U+63B4 <cjk>
	0xCE: [`\u69FB`].string() // U+69FB <cjk>
	0xCF: [`\u4F43`].string() // U+4F43 <cjk>
	0xD0: [`\u6F2C`].string() // U+6F2C <cjk>
	0xD1: [`\u67D8`].string() // U+67D8 <cjk>
	0xD2: [`\u8FBB`].string() // U+8FBB <cjk>
	0xD3: [`\u8526`].string() // U+8526 <cjk>
	0xD4: [`\u7DB4`].string() // U+7DB4 <cjk>
	0xD5: [`\u9354`].string() // U+9354 <cjk>
	0xD6: [`\u693F`].string() // U+693F <cjk>
	0xD7: [`\u6F70`].string() // U+6F70 <cjk>
	0xD8: [`\u576A`].string() // U+576A <cjk>
	0xD9: [`\u58F7`].string() // U+58F7 <cjk>
	0xDA: [`\u5B2C`].string() // U+5B2C <cjk>
	0xDB: [`\u7D2C`].string() // U+7D2C <cjk>
	0xDC: [`\u722A`].string() // U+722A <cjk>
	0xDD: [`\u540A`].string() // U+540A <cjk>
	0xDE: [`\u91E3`].string() // U+91E3 <cjk>
	0xDF: [`\u9DB4`].string() // U+9DB4 <cjk>
	0xE0: [`\u4EAD`].string() // U+4EAD <cjk>
	0xE1: [`\u4F4E`].string() // U+4F4E <cjk>
	0xE2: [`\u505C`].string() // U+505C <cjk>
	0xE3: [`\u5075`].string() // U+5075 <cjk>
	0xE4: [`\u5243`].string() // U+5243 <cjk>
	0xE5: [`\u8C9E`].string() // U+8C9E <cjk>
	0xE6: [`\u5448`].string() // U+5448 <cjk>
	0xE7: [`\u5824`].string() // U+5824 <cjk>
	0xE8: [`\u5B9A`].string() // U+5B9A <cjk>
	0xE9: [`\u5E1D`].string() // U+5E1D <cjk>
	0xEA: [`\u5E95`].string() // U+5E95 <cjk>
	0xEB: [`\u5EAD`].string() // U+5EAD <cjk>
	0xEC: [`\u5EF7`].string() // U+5EF7 <cjk>
	0xED: [`\u5F1F`].string() // U+5F1F <cjk>
	0xEE: [`\u608C`].string() // U+608C <cjk>
	0xEF: [`\u62B5`].string() // U+62B5 <cjk>
	0xF0: [`\u633A`].string() // U+633A <cjk>
	0xF1: [`\u63D0`].string() // U+63D0 <cjk>
	0xF2: [`\u68AF`].string() // U+68AF <cjk>
	0xF3: [`\u6C40`].string() // U+6C40 <cjk>
	0xF4: [`\u7887`].string() // U+7887 <cjk>
	0xF5: [`\u798E`].string() // U+798E <cjk>
	0xF6: [`\u7A0B`].string() // U+7A0B <cjk>
	0xF7: [`\u7DE0`].string() // U+7DE0 <cjk>
	0xF8: [`\u8247`].string() // U+8247 <cjk>
	0xF9: [`\u8A02`].string() // U+8A02 <cjk>
	0xFA: [`\u8AE6`].string() // U+8AE6 <cjk>
	0xFB: [`\u8E44`].string() // U+8E44 <cjk>
	0xFC: [`\u9013`].string() // U+9013 <cjk>
}

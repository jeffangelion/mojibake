module mojibake

const jis_x_0213_doublebyte_0x82 = {
	0x40: [`\u25B7`].string() // U+25B7 WHITE RIGHT-POINTING TRIANGLE
	0x41: [`\u25B6`].string() // U+25B6 BLACK RIGHT-POINTING TRIANGLE
	0x42: [`\u25C1`].string() // U+25C1 WHITE LEFT-POINTING TRIANGLE
	0x43: [`\u25C0`].string() // U+25C0 BLACK LEFT-POINTING TRIANGLE
	0x44: [`\u2197`].string() // U+2197 NORTH EAST ARROW
	0x45: [`\u2198`].string() // U+2198 SOUTH EAST ARROW
	0x46: [`\u2196`].string() // U+2196 NORTH WEST ARROW
	0x47: [`\u2199`].string() // U+2199 SOUTH WEST ARROW
	0x48: [`\u21C4`].string() // U+21C4 RIGHTWARDS ARROW OVER LEFTWARDS ARROW
	0x49: [`\u21E8`].string() // U+21E8 RIGHTWARDS WHITE ARROW
	0x4A: [`\u21E6`].string() // U+21E6 LEFTWARDS WHITE ARROW
	0x4B: [`\u21E7`].string() // U+21E7 UPWARDS WHITE ARROW
	0x4C: [`\u21E9`].string() // U+21E9 DOWNWARDS WHITE ARROW
	0x4D: [`\u2934`].string() // U+2934 ARROW POINTING RIGHTWARDS THEN CURVING UPWARDS
	0x4E: [`\u2935`].string() // U+2935 ARROW POINTING RIGHTWARDS THEN CURVING DOWNWARDS
	0x4F: [`\uFF10`].string() // U+FF10 FULLWIDTH DIGIT ZERO
	0x50: [`\uFF11`].string() // U+FF11 FULLWIDTH DIGIT ONE
	0x51: [`\uFF12`].string() // U+FF12 FULLWIDTH DIGIT TWO
	0x52: [`\uFF13`].string() // U+FF13 FULLWIDTH DIGIT THREE
	0x53: [`\uFF14`].string() // U+FF14 FULLWIDTH DIGIT FOUR
	0x54: [`\uFF15`].string() // U+FF15 FULLWIDTH DIGIT FIVE
	0x55: [`\uFF16`].string() // U+FF16 FULLWIDTH DIGIT SIX
	0x56: [`\uFF17`].string() // U+FF17 FULLWIDTH DIGIT SEVEN
	0x57: [`\uFF18`].string() // U+FF18 FULLWIDTH DIGIT EIGHT
	0x58: [`\uFF19`].string() // U+FF19 FULLWIDTH DIGIT NINE
	0x59: [`\u29BF`].string() // U+29BF CIRCLED BULLET
	0x5A: [`\u25C9`].string() // U+25C9 FISHEYE
	0x5B: [`\u303D`].string() // U+303D PART ALTERNATION MARK
	0x5C: [`\uFE46`].string() // U+FE46 WHITE SESAME DOT
	0x5D: [`\uFE45`].string() // U+FE45 SESAME DOT
	0x5E: [`\u25E6`].string() // U+25E6 WHITE BULLET
	0x5F: [`\u2022`].string() // U+2022 BULLET
	0x60: [`\uFF21`].string() // U+FF21 FULLWIDTH LATIN CAPITAL LETTER A
	0x61: [`\uFF22`].string() // U+FF22 FULLWIDTH LATIN CAPITAL LETTER B
	0x62: [`\uFF23`].string() // U+FF23 FULLWIDTH LATIN CAPITAL LETTER C
	0x63: [`\uFF24`].string() // U+FF24 FULLWIDTH LATIN CAPITAL LETTER D
	0x64: [`\uFF25`].string() // U+FF25 FULLWIDTH LATIN CAPITAL LETTER E
	0x65: [`\uFF26`].string() // U+FF26 FULLWIDTH LATIN CAPITAL LETTER F
	0x66: [`\uFF27`].string() // U+FF27 FULLWIDTH LATIN CAPITAL LETTER G
	0x67: [`\uFF28`].string() // U+FF28 FULLWIDTH LATIN CAPITAL LETTER H
	0x68: [`\uFF29`].string() // U+FF29 FULLWIDTH LATIN CAPITAL LETTER I
	0x69: [`\uFF2A`].string() // U+FF2A FULLWIDTH LATIN CAPITAL LETTER J
	0x6A: [`\uFF2B`].string() // U+FF2B FULLWIDTH LATIN CAPITAL LETTER K
	0x6B: [`\uFF2C`].string() // U+FF2C FULLWIDTH LATIN CAPITAL LETTER L
	0x6C: [`\uFF2D`].string() // U+FF2D FULLWIDTH LATIN CAPITAL LETTER M
	0x6D: [`\uFF2E`].string() // U+FF2E FULLWIDTH LATIN CAPITAL LETTER N
	0x6E: [`\uFF2F`].string() // U+FF2F FULLWIDTH LATIN CAPITAL LETTER O
	0x6F: [`\uFF30`].string() // U+FF30 FULLWIDTH LATIN CAPITAL LETTER P
	0x70: [`\uFF31`].string() // U+FF31 FULLWIDTH LATIN CAPITAL LETTER Q
	0x71: [`\uFF32`].string() // U+FF32 FULLWIDTH LATIN CAPITAL LETTER R
	0x72: [`\uFF33`].string() // U+FF33 FULLWIDTH LATIN CAPITAL LETTER S
	0x73: [`\uFF34`].string() // U+FF34 FULLWIDTH LATIN CAPITAL LETTER T
	0x74: [`\uFF35`].string() // U+FF35 FULLWIDTH LATIN CAPITAL LETTER U
	0x75: [`\uFF36`].string() // U+FF36 FULLWIDTH LATIN CAPITAL LETTER V
	0x76: [`\uFF37`].string() // U+FF37 FULLWIDTH LATIN CAPITAL LETTER W
	0x77: [`\uFF38`].string() // U+FF38 FULLWIDTH LATIN CAPITAL LETTER X
	0x78: [`\uFF39`].string() // U+FF39 FULLWIDTH LATIN CAPITAL LETTER Y
	0x79: [`\uFF3A`].string() // U+FF3A FULLWIDTH LATIN CAPITAL LETTER Z
	0x7A: [`\u2213`].string() // U+2213 MINUS-OR-PLUS SIGN
	0x7B: [`\u2135`].string() // U+2135 ALEF SYMBOL
	0x7C: [`\u210F`].string() // U+210F PLANCK CONSTANT OVER TWO PI
	0x7D: [`\u33CB`].string() // U+33CB SQUARE HP
	0x7E: [`\u2113`].string() // U+2113 SCRIPT SMALL L
	0x80: [`\u2127`].string() // U+2127 INVERTED OHM SIGN
	0x81: [`\uFF41`].string() // U+FF41 FULLWIDTH LATIN SMALL LETTER A
	0x82: [`\uFF42`].string() // U+FF42 FULLWIDTH LATIN SMALL LETTER B
	0x83: [`\uFF43`].string() // U+FF43 FULLWIDTH LATIN SMALL LETTER C
	0x84: [`\uFF44`].string() // U+FF44 FULLWIDTH LATIN SMALL LETTER D
	0x85: [`\uFF45`].string() // U+FF45 FULLWIDTH LATIN SMALL LETTER E
	0x86: [`\uFF46`].string() // U+FF46 FULLWIDTH LATIN SMALL LETTER F
	0x87: [`\uFF47`].string() // U+FF47 FULLWIDTH LATIN SMALL LETTER G
	0x88: [`\uFF48`].string() // U+FF48 FULLWIDTH LATIN SMALL LETTER H
	0x89: [`\uFF49`].string() // U+FF49 FULLWIDTH LATIN SMALL LETTER I
	0x8A: [`\uFF4A`].string() // U+FF4A FULLWIDTH LATIN SMALL LETTER J
	0x8B: [`\uFF4B`].string() // U+FF4B FULLWIDTH LATIN SMALL LETTER K
	0x8C: [`\uFF4C`].string() // U+FF4C FULLWIDTH LATIN SMALL LETTER L
	0x8D: [`\uFF4D`].string() // U+FF4D FULLWIDTH LATIN SMALL LETTER M
	0x8E: [`\uFF4E`].string() // U+FF4E FULLWIDTH LATIN SMALL LETTER N
	0x8F: [`\uFF4F`].string() // U+FF4F FULLWIDTH LATIN SMALL LETTER O
	0x90: [`\uFF50`].string() // U+FF50 FULLWIDTH LATIN SMALL LETTER P
	0x91: [`\uFF51`].string() // U+FF51 FULLWIDTH LATIN SMALL LETTER Q
	0x92: [`\uFF52`].string() // U+FF52 FULLWIDTH LATIN SMALL LETTER R
	0x93: [`\uFF53`].string() // U+FF53 FULLWIDTH LATIN SMALL LETTER S
	0x94: [`\uFF54`].string() // U+FF54 FULLWIDTH LATIN SMALL LETTER T
	0x95: [`\uFF55`].string() // U+FF55 FULLWIDTH LATIN SMALL LETTER U
	0x96: [`\uFF56`].string() // U+FF56 FULLWIDTH LATIN SMALL LETTER V
	0x97: [`\uFF57`].string() // U+FF57 FULLWIDTH LATIN SMALL LETTER W
	0x98: [`\uFF58`].string() // U+FF58 FULLWIDTH LATIN SMALL LETTER X
	0x99: [`\uFF59`].string() // U+FF59 FULLWIDTH LATIN SMALL LETTER Y
	0x9A: [`\uFF5A`].string() // U+FF5A FULLWIDTH LATIN SMALL LETTER Z
	0x9B: [`\u30A0`].string() // U+30A0 KATAKANA-HIRAGANA DOUBLE HYPHEN
	0x9C: [`\u2013`].string() // U+2013 EN DASH
	0x9D: [`\u29FA`].string() // U+29FA DOUBLE PLUS
	0x9E: [`\u29FB`].string() // U+29FB TRIPLE PLUS
	0x9F: [`\u3041`].string() // U+3041 HIRAGANA LETTER SMALL A
	0xA0: [`\u3042`].string() // U+3042 HIRAGANA LETTER A
	0xA1: [`\u3043`].string() // U+3043 HIRAGANA LETTER SMALL I
	0xA2: [`\u3044`].string() // U+3044 HIRAGANA LETTER I
	0xA3: [`\u3045`].string() // U+3045 HIRAGANA LETTER SMALL U
	0xA4: [`\u3046`].string() // U+3046 HIRAGANA LETTER U
	0xA5: [`\u3047`].string() // U+3047 HIRAGANA LETTER SMALL E
	0xA6: [`\u3048`].string() // U+3048 HIRAGANA LETTER E
	0xA7: [`\u3049`].string() // U+3049 HIRAGANA LETTER SMALL O
	0xA8: [`\u304A`].string() // U+304A HIRAGANA LETTER O
	0xA9: [`\u304B`].string() // U+304B HIRAGANA LETTER KA
	0xAA: [`\u304C`].string() // U+304C HIRAGANA LETTER GA
	0xAB: [`\u304D`].string() // U+304D HIRAGANA LETTER KI
	0xAC: [`\u304E`].string() // U+304E HIRAGANA LETTER GI
	0xAD: [`\u304F`].string() // U+304F HIRAGANA LETTER KU
	0xAE: [`\u3050`].string() // U+3050 HIRAGANA LETTER GU
	0xAF: [`\u3051`].string() // U+3051 HIRAGANA LETTER KE
	0xB0: [`\u3052`].string() // U+3052 HIRAGANA LETTER GE
	0xB1: [`\u3053`].string() // U+3053 HIRAGANA LETTER KO
	0xB2: [`\u3054`].string() // U+3054 HIRAGANA LETTER GO
	0xB3: [`\u3055`].string() // U+3055 HIRAGANA LETTER SA
	0xB4: [`\u3056`].string() // U+3056 HIRAGANA LETTER ZA
	0xB5: [`\u3057`].string() // U+3057 HIRAGANA LETTER SI
	0xB6: [`\u3058`].string() // U+3058 HIRAGANA LETTER ZI
	0xB7: [`\u3059`].string() // U+3059 HIRAGANA LETTER SU
	0xB8: [`\u305A`].string() // U+305A HIRAGANA LETTER ZU
	0xB9: [`\u305B`].string() // U+305B HIRAGANA LETTER SE
	0xBA: [`\u305C`].string() // U+305C HIRAGANA LETTER ZE
	0xBB: [`\u305D`].string() // U+305D HIRAGANA LETTER SO
	0xBC: [`\u305E`].string() // U+305E HIRAGANA LETTER ZO
	0xBD: [`\u305F`].string() // U+305F HIRAGANA LETTER TA
	0xBE: [`\u3060`].string() // U+3060 HIRAGANA LETTER DA
	0xBF: [`\u3061`].string() // U+3061 HIRAGANA LETTER TI
	0xC0: [`\u3062`].string() // U+3062 HIRAGANA LETTER DI
	0xC1: [`\u3063`].string() // U+3063 HIRAGANA LETTER SMALL TU
	0xC2: [`\u3064`].string() // U+3064 HIRAGANA LETTER TU
	0xC3: [`\u3065`].string() // U+3065 HIRAGANA LETTER DU
	0xC4: [`\u3066`].string() // U+3066 HIRAGANA LETTER TE
	0xC5: [`\u3067`].string() // U+3067 HIRAGANA LETTER DE
	0xC6: [`\u3068`].string() // U+3068 HIRAGANA LETTER TO
	0xC7: [`\u3069`].string() // U+3069 HIRAGANA LETTER DO
	0xC8: [`\u306A`].string() // U+306A HIRAGANA LETTER NA
	0xC9: [`\u306B`].string() // U+306B HIRAGANA LETTER NI
	0xCA: [`\u306C`].string() // U+306C HIRAGANA LETTER NU
	0xCB: [`\u306D`].string() // U+306D HIRAGANA LETTER NE
	0xCC: [`\u306E`].string() // U+306E HIRAGANA LETTER NO
	0xCD: [`\u306F`].string() // U+306F HIRAGANA LETTER HA
	0xCE: [`\u3070`].string() // U+3070 HIRAGANA LETTER BA
	0xCF: [`\u3071`].string() // U+3071 HIRAGANA LETTER PA
	0xD0: [`\u3072`].string() // U+3072 HIRAGANA LETTER HI
	0xD1: [`\u3073`].string() // U+3073 HIRAGANA LETTER BI
	0xD2: [`\u3074`].string() // U+3074 HIRAGANA LETTER PI
	0xD3: [`\u3075`].string() // U+3075 HIRAGANA LETTER HU
	0xD4: [`\u3076`].string() // U+3076 HIRAGANA LETTER BU
	0xD5: [`\u3077`].string() // U+3077 HIRAGANA LETTER PU
	0xD6: [`\u3078`].string() // U+3078 HIRAGANA LETTER HE
	0xD7: [`\u3079`].string() // U+3079 HIRAGANA LETTER BE
	0xD8: [`\u307A`].string() // U+307A HIRAGANA LETTER PE
	0xD9: [`\u307B`].string() // U+307B HIRAGANA LETTER HO
	0xDA: [`\u307C`].string() // U+307C HIRAGANA LETTER BO
	0xDB: [`\u307D`].string() // U+307D HIRAGANA LETTER PO
	0xDC: [`\u307E`].string() // U+307E HIRAGANA LETTER MA
	0xDD: [`\u307F`].string() // U+307F HIRAGANA LETTER MI
	0xDE: [`\u3080`].string() // U+3080 HIRAGANA LETTER MU
	0xDF: [`\u3081`].string() // U+3081 HIRAGANA LETTER ME
	0xE0: [`\u3082`].string() // U+3082 HIRAGANA LETTER MO
	0xE1: [`\u3083`].string() // U+3083 HIRAGANA LETTER SMALL YA
	0xE2: [`\u3084`].string() // U+3084 HIRAGANA LETTER YA
	0xE3: [`\u3085`].string() // U+3085 HIRAGANA LETTER SMALL YU
	0xE4: [`\u3086`].string() // U+3086 HIRAGANA LETTER YU
	0xE5: [`\u3087`].string() // U+3087 HIRAGANA LETTER SMALL YO
	0xE6: [`\u3088`].string() // U+3088 HIRAGANA LETTER YO
	0xE7: [`\u3089`].string() // U+3089 HIRAGANA LETTER RA
	0xE8: [`\u308A`].string() // U+308A HIRAGANA LETTER RI
	0xE9: [`\u308B`].string() // U+308B HIRAGANA LETTER RU
	0xEA: [`\u308C`].string() // U+308C HIRAGANA LETTER RE
	0xEB: [`\u308D`].string() // U+308D HIRAGANA LETTER RO
	0xEC: [`\u308E`].string() // U+308E HIRAGANA LETTER SMALL WA
	0xED: [`\u308F`].string() // U+308F HIRAGANA LETTER WA
	0xEE: [`\u3090`].string() // U+3090 HIRAGANA LETTER WI
	0xEF: [`\u3091`].string() // U+3091 HIRAGANA LETTER WE
	0xF0: [`\u3092`].string() // U+3092 HIRAGANA LETTER WO
	0xF1: [`\u3093`].string() // U+3093 HIRAGANA LETTER N
	0xF2: [`\u3094`].string() // U+3094 HIRAGANA LETTER VU
	0xF3: [`\u3095`].string() // U+3095 HIRAGANA LETTER SMALL KA
	0xF4: [`\u3096`].string() // U+3096 HIRAGANA LETTER SMALL KE
	0xF5: [`\u304B`,`\u309A`].string() // U+304B+309A
	0xF6: [`\u304D`,`\u309A`].string() // U+304D+309A
	0xF7: [`\u304F`,`\u309A`].string() // U+304F+309A
	0xF8: [`\u3051`,`\u309A`].string() // U+3051+309A
	0xF9: [`\u3053`,`\u309A`].string() // U+3053+309A
}

module mojibake

const jis_x_0213_doublebyte_0xef = {
	0x40: [`\u91E5`].string() // U+91E5 <cjk>
	0x41: [`\u91ED`].string() // U+91ED <cjk>
	0x42: [`\u91F1`].string() // U+91F1 <cjk>
	0x43: [`\u9207`].string() // U+9207 <cjk>
	0x44: [`\u9210`].string() // U+9210 <cjk>
	0x45: [`\u9238`].string() // U+9238 <cjk>
	0x46: [`\u9239`].string() // U+9239 <cjk>
	0x47: [`\u923A`].string() // U+923A <cjk>
	0x48: [`\u923C`].string() // U+923C <cjk>
	0x49: [`\u9240`].string() // U+9240 <cjk>
	0x4A: [`\u9243`].string() // U+9243 <cjk>
	0x4B: [`\u924F`].string() // U+924F <cjk>
	0x4C: [`\u9278`].string() // U+9278 <cjk>
	0x4D: [`\u9288`].string() // U+9288 <cjk>
	0x4E: [`\u92C2`].string() // U+92C2 <cjk>
	0x4F: [`\u92CB`].string() // U+92CB <cjk>
	0x50: [`\u92CC`].string() // U+92CC <cjk>
	0x51: [`\u92D3`].string() // U+92D3 <cjk>
	0x52: [`\u92E0`].string() // U+92E0 <cjk>
	0x53: [`\u92FF`].string() // U+92FF <cjk>
	0x54: [`\u9304`].string() // U+9304 <cjk>
	0x55: [`\u931F`].string() // U+931F <cjk>
	0x56: [`\u9321`].string() // U+9321 <cjk>
	0x57: [`\u9325`].string() // U+9325 <cjk>
	0x58: [`\u9348`].string() // U+9348 <cjk>
	0x59: [`\u9349`].string() // U+9349 <cjk>
	0x5A: [`\u934A`].string() // U+934A <cjk>
	0x5B: [`\u9364`].string() // U+9364 <cjk>
	0x5C: [`\u9365`].string() // U+9365 <cjk>
	0x5D: [`\u936A`].string() // U+936A <cjk>
	0x5E: [`\u9370`].string() // U+9370 <cjk>
	0x5F: [`\u939B`].string() // U+939B <cjk>
	0x60: [`\u93A3`].string() // U+93A3 <cjk>
	0x61: [`\u93BA`].string() // U+93BA <cjk>
	0x62: [`\u93C6`].string() // U+93C6 <cjk>
	0x63: [`\u93DE`].string() // U+93DE <cjk>
	0x64: [`\u93DF`].string() // U+93DF <cjk>
	0x65: [`\u9404`].string() // U+9404 <cjk>
	0x66: [`\u93FD`].string() // U+93FD <cjk>
	0x67: [`\u9433`].string() // U+9433 <cjk>
	0x68: [`\u944A`].string() // U+944A <cjk>
	0x69: [`\u9463`].string() // U+9463 <cjk>
	0x6A: [`\u946B`].string() // U+946B <cjk>
	0x6B: [`\u9471`].string() // U+9471 <cjk>
	0x6C: [`\u9472`].string() // U+9472 <cjk>
	0x6D: [`\u958E`].string() // U+958E <cjk>
	0x6E: [`\u959F`].string() // U+959F <cjk>
	0x6F: [`\u95A6`].string() // U+95A6 <cjk>
	0x70: [`\u95A9`].string() // U+95A9 <cjk>
	0x71: [`\u95AC`].string() // U+95AC <cjk>
	0x72: [`\u95B6`].string() // U+95B6 <cjk>
	0x73: [`\u95BD`].string() // U+95BD <cjk>
	0x74: [`\u95CB`].string() // U+95CB <cjk>
	0x75: [`\u95D0`].string() // U+95D0 <cjk>
	0x76: [`\u95D3`].string() // U+95D3 <cjk>
	0x77: [`\u49B0`].string() // U+49B0 <cjk>
	0x78: [`\u95DA`].string() // U+95DA <cjk>
	0x79: [`\u95DE`].string() // U+95DE <cjk>
	0x7A: [`\u9658`].string() // U+9658 <cjk>
	0x7B: [`\u9684`].string() // U+9684 <cjk>
	0x7C: [`\uF9DC`].string() // U+F9DC CJK COMPATIBILITY IDEOGRAPH-F9DC
	0x7D: [`\u969D`].string() // U+969D <cjk>
	0x7E: [`\u96A4`].string() // U+96A4 <cjk>
	0x80: [`\u96A5`].string() // U+96A5 <cjk>
	0x81: [`\u96D2`].string() // U+96D2 <cjk>
	0x82: [`\u96DE`].string() // U+96DE <cjk>
	0x83: [`\uFA68`].string() // U+FA68 CJK COMPATIBILITY IDEOGRAPH-FA68
	0x84: [`\u96E9`].string() // U+96E9 <cjk>
	0x85: [`\u96EF`].string() // U+96EF <cjk>
	0x86: [`\u9733`].string() // U+9733 <cjk>
	0x87: [`\u973B`].string() // U+973B <cjk>
	0x88: [`\u974D`].string() // U+974D <cjk>
	0x89: [`\u974E`].string() // U+974E <cjk>
	0x8A: [`\u974F`].string() // U+974F <cjk>
	0x8B: [`\u975A`].string() // U+975A <cjk>
	0x8C: [`\u976E`].string() // U+976E <cjk>
	0x8D: [`\u9773`].string() // U+9773 <cjk>
	0x8E: [`\u9795`].string() // U+9795 <cjk>
	0x8F: [`\u97AE`].string() // U+97AE <cjk>
	0x90: [`\u97BA`].string() // U+97BA <cjk>
	0x91: [`\u97C1`].string() // U+97C1 <cjk>
	0x92: [`\u97C9`].string() // U+97C9 <cjk>
	0x93: [`\u97DE`].string() // U+97DE <cjk>
	0x94: [`\u97DB`].string() // U+97DB <cjk>
	0x95: [`\u97F4`].string() // U+97F4 <cjk>
	0x96: [`\uFA69`].string() // U+FA69 CJK COMPATIBILITY IDEOGRAPH-FA69
	0x97: [`\u980A`].string() // U+980A <cjk>
	0x98: [`\u981E`].string() // U+981E <cjk>
	0x99: [`\u982B`].string() // U+982B <cjk>
	0x9A: [`\u9830`].string() // U+9830 <cjk>
	0x9B: [`\uFA6A`].string() // U+FA6A CJK COMPATIBILITY IDEOGRAPH-FA6A
	0x9C: [`\u9852`].string() // U+9852 <cjk>
	0x9D: [`\u9853`].string() // U+9853 <cjk>
	0x9E: [`\u9856`].string() // U+9856 <cjk>
	0x9F: [`\u9857`].string() // U+9857 <cjk>
	0xA0: [`\u9859`].string() // U+9859 <cjk>
	0xA1: [`\u985A`].string() // U+985A <cjk>
	0xA2: [`\uF9D0`].string() // U+F9D0 CJK COMPATIBILITY IDEOGRAPH-F9D0
	0xA3: [`\u9865`].string() // U+9865 <cjk>
	0xA4: [`\u986C`].string() // U+986C <cjk>
	0xA5: [`\u98BA`].string() // U+98BA <cjk>
	0xA6: [`\u98C8`].string() // U+98C8 <cjk>
	0xA7: [`\u98E7`].string() // U+98E7 <cjk>
	0xA8: [`\u9958`].string() // U+9958 <cjk>
	0xA9: [`\u999E`].string() // U+999E <cjk>
	0xAA: [`\u9A02`].string() // U+9A02 <cjk>
	0xAB: [`\u9A03`].string() // U+9A03 <cjk>
	0xAC: [`\u9A24`].string() // U+9A24 <cjk>
	0xAD: [`\u9A2D`].string() // U+9A2D <cjk>
	0xAE: [`\u9A2E`].string() // U+9A2E <cjk>
	0xAF: [`\u9A38`].string() // U+9A38 <cjk>
	0xB0: [`\u9A4A`].string() // U+9A4A <cjk>
	0xB1: [`\u9A4E`].string() // U+9A4E <cjk>
	0xB2: [`\u9A52`].string() // U+9A52 <cjk>
	0xB3: [`\u9AB6`].string() // U+9AB6 <cjk>
	0xB4: [`\u9AC1`].string() // U+9AC1 <cjk>
	0xB5: [`\u9AC3`].string() // U+9AC3 <cjk>
	0xB6: [`\u9ACE`].string() // U+9ACE <cjk>
	0xB7: [`\u9AD6`].string() // U+9AD6 <cjk>
	0xB8: [`\u9AF9`].string() // U+9AF9 <cjk>
	0xB9: [`\u9B02`].string() // U+9B02 <cjk>
	0xBA: [`\u9B08`].string() // U+9B08 <cjk>
	0xBB: [`\u9B20`].string() // U+9B20 <cjk>
	0xBC: [`\u4C17`].string() // U+4C17 <cjk>
	0xBD: [`\u9B2D`].string() // U+9B2D <cjk>
	0xBE: [`\u9B5E`].string() // U+9B5E <cjk>
	0xBF: [`\u9B79`].string() // U+9B79 <cjk>
	0xC0: [`\u9B66`].string() // U+9B66 <cjk>
	0xC1: [`\u9B72`].string() // U+9B72 <cjk>
	0xC2: [`\u9B75`].string() // U+9B75 <cjk>
	0xC3: [`\u9B84`].string() // U+9B84 <cjk>
	0xC4: [`\u9B8A`].string() // U+9B8A <cjk>
	0xC5: [`\u9B8F`].string() // U+9B8F <cjk>
	0xC6: [`\u9B9E`].string() // U+9B9E <cjk>
	0xC7: [`\u9BA7`].string() // U+9BA7 <cjk>
	0xC8: [`\u9BC1`].string() // U+9BC1 <cjk>
	0xC9: [`\u9BCE`].string() // U+9BCE <cjk>
	0xCA: [`\u9BE5`].string() // U+9BE5 <cjk>
	0xCB: [`\u9BF8`].string() // U+9BF8 <cjk>
	0xCC: [`\u9BFD`].string() // U+9BFD <cjk>
	0xCD: [`\u9C00`].string() // U+9C00 <cjk>
	0xCE: [`\u9C23`].string() // U+9C23 <cjk>
	0xCF: [`\u9C41`].string() // U+9C41 <cjk>
	0xD0: [`\u9C4F`].string() // U+9C4F <cjk>
	0xD1: [`\u9C50`].string() // U+9C50 <cjk>
	0xD2: [`\u9C53`].string() // U+9C53 <cjk>
	0xD3: [`\u9C63`].string() // U+9C63 <cjk>
	0xD4: [`\u9C65`].string() // U+9C65 <cjk>
	0xD5: [`\u9C77`].string() // U+9C77 <cjk>
	0xD6: [`\u9D1D`].string() // U+9D1D <cjk>
	0xD7: [`\u9D1E`].string() // U+9D1E <cjk>
	0xD8: [`\u9D43`].string() // U+9D43 <cjk>
	0xD9: [`\u9D47`].string() // U+9D47 <cjk>
	0xDA: [`\u9D52`].string() // U+9D52 <cjk>
	0xDB: [`\u9D63`].string() // U+9D63 <cjk>
	0xDC: [`\u9D70`].string() // U+9D70 <cjk>
	0xDD: [`\u9D7C`].string() // U+9D7C <cjk>
	0xDE: [`\u9D8A`].string() // U+9D8A <cjk>
	0xDF: [`\u9D96`].string() // U+9D96 <cjk>
	0xE0: [`\u9DC0`].string() // U+9DC0 <cjk>
	0xE1: [`\u9DAC`].string() // U+9DAC <cjk>
	0xE2: [`\u9DBC`].string() // U+9DBC <cjk>
	0xE3: [`\u9DD7`].string() // U+9DD7 <cjk>
	0xE4: utf32_to_str(0x2A190) // U+2A190 <cjk>
	0xE5: [`\u9DE7`].string() // U+9DE7 <cjk>
	0xE6: [`\u9E07`].string() // U+9E07 <cjk>
	0xE7: [`\u9E15`].string() // U+9E15 <cjk>
	0xE8: [`\u9E7C`].string() // U+9E7C <cjk>
	0xE9: [`\u9E9E`].string() // U+9E9E <cjk>
	0xEA: [`\u9EA4`].string() // U+9EA4 <cjk>
	0xEB: [`\u9EAC`].string() // U+9EAC <cjk>
	0xEC: [`\u9EAF`].string() // U+9EAF <cjk>
	0xED: [`\u9EB4`].string() // U+9EB4 <cjk>
	0xEE: [`\u9EB5`].string() // U+9EB5 <cjk>
	0xEF: [`\u9EC3`].string() // U+9EC3 <cjk>
	0xF0: [`\u9ED1`].string() // U+9ED1 <cjk>
	0xF1: [`\u9F10`].string() // U+9F10 <cjk>
	0xF2: [`\u9F39`].string() // U+9F39 <cjk>
	0xF3: [`\u9F57`].string() // U+9F57 <cjk>
	0xF4: [`\u9F90`].string() // U+9F90 <cjk>
	0xF5: [`\u9F94`].string() // U+9F94 <cjk>
	0xF6: [`\u9F97`].string() // U+9F97 <cjk>
	0xF7: [`\u9FA2`].string() // U+9FA2 <cjk>
	0xF8: [`\u59F8`].string() // U+59F8 <cjk>
	0xF9: [`\u5C5B`].string() // U+5C5B <cjk>
	0xFA: [`\u5E77`].string() // U+5E77 <cjk>
	0xFB: [`\u7626`].string() // U+7626 <cjk>
	0xFC: [`\u7E6B`].string() // U+7E6B <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xf6 = {
	0x40: [`\u74A0`].string() // U+74A0 <cjk>
	0x41: [`\u74A1`].string() // U+74A1 <cjk>
	0x42: [`\u74A5`].string() // U+74A5 <cjk>
	0x43: [`\u74AA`].string() // U+74AA <cjk>
	0x44: [`\u74AB`].string() // U+74AB <cjk>
	0x45: [`\u74B9`].string() // U+74B9 <cjk>
	0x46: [`\u74BB`].string() // U+74BB <cjk>
	0x47: [`\u74BA`].string() // U+74BA <cjk>
	0x48: [`\u74D6`].string() // U+74D6 <cjk>
	0x49: [`\u74D8`].string() // U+74D8 <cjk>
	0x4A: [`\u74DE`].string() // U+74DE <cjk>
	0x4B: [`\u74EF`].string() // U+74EF <cjk>
	0x4C: [`\u74EB`].string() // U+74EB <cjk>
	0x4D: utf32_to_str(0x24B56) // U+24B56 <cjk>
	0x4E: [`\u74FA`].string() // U+74FA <cjk>
	0x4F: utf32_to_str(0x24B6F) // U+24B6F <cjk>
	0x50: [`\u7520`].string() // U+7520 <cjk>
	0x51: [`\u7524`].string() // U+7524 <cjk>
	0x52: [`\u752A`].string() // U+752A <cjk>
	0x53: [`\u3F57`].string() // U+3F57 <cjk>
	0x54: utf32_to_str(0x24C16) // U+24C16 <cjk>
	0x55: [`\u753D`].string() // U+753D <cjk>
	0x56: [`\u753E`].string() // U+753E <cjk>
	0x57: [`\u7540`].string() // U+7540 <cjk>
	0x58: [`\u7548`].string() // U+7548 <cjk>
	0x59: [`\u754E`].string() // U+754E <cjk>
	0x5A: [`\u7550`].string() // U+7550 <cjk>
	0x5B: [`\u7552`].string() // U+7552 <cjk>
	0x5C: [`\u756C`].string() // U+756C <cjk>
	0x5D: [`\u7572`].string() // U+7572 <cjk>
	0x5E: [`\u7571`].string() // U+7571 <cjk>
	0x5F: [`\u757A`].string() // U+757A <cjk>
	0x60: [`\u757D`].string() // U+757D <cjk>
	0x61: [`\u757E`].string() // U+757E <cjk>
	0x62: [`\u7581`].string() // U+7581 <cjk>
	0x63: utf32_to_str(0x24D14) // U+24D14 <cjk>
	0x64: [`\u758C`].string() // U+758C <cjk>
	0x65: [`\u3F75`].string() // U+3F75 <cjk>
	0x66: [`\u75A2`].string() // U+75A2 <cjk>
	0x67: [`\u3F77`].string() // U+3F77 <cjk>
	0x68: [`\u75B0`].string() // U+75B0 <cjk>
	0x69: [`\u75B7`].string() // U+75B7 <cjk>
	0x6A: [`\u75BF`].string() // U+75BF <cjk>
	0x6B: [`\u75C0`].string() // U+75C0 <cjk>
	0x6C: [`\u75C6`].string() // U+75C6 <cjk>
	0x6D: [`\u75CF`].string() // U+75CF <cjk>
	0x6E: [`\u75D3`].string() // U+75D3 <cjk>
	0x6F: [`\u75DD`].string() // U+75DD <cjk>
	0x70: [`\u75DF`].string() // U+75DF <cjk>
	0x71: [`\u75E0`].string() // U+75E0 <cjk>
	0x72: [`\u75E7`].string() // U+75E7 <cjk>
	0x73: [`\u75EC`].string() // U+75EC <cjk>
	0x74: [`\u75EE`].string() // U+75EE <cjk>
	0x75: [`\u75F1`].string() // U+75F1 <cjk>
	0x76: [`\u75F9`].string() // U+75F9 <cjk>
	0x77: [`\u7603`].string() // U+7603 <cjk>
	0x78: [`\u7618`].string() // U+7618 <cjk>
	0x79: [`\u7607`].string() // U+7607 <cjk>
	0x7A: [`\u760F`].string() // U+760F <cjk>
	0x7B: [`\u3FAE`].string() // U+3FAE <cjk>
	0x7C: utf32_to_str(0x24E0E) // U+24E0E <cjk>
	0x7D: [`\u7613`].string() // U+7613 <cjk>
	0x7E: [`\u761B`].string() // U+761B <cjk>
	0x80: [`\u761C`].string() // U+761C <cjk>
	0x81: utf32_to_str(0x24E37) // U+24E37 <cjk>
	0x82: [`\u7625`].string() // U+7625 <cjk>
	0x83: [`\u7628`].string() // U+7628 <cjk>
	0x84: [`\u763C`].string() // U+763C <cjk>
	0x85: [`\u7633`].string() // U+7633 <cjk>
	0x86: utf32_to_str(0x24E6A) // U+24E6A <cjk>
	0x87: [`\u3FC9`].string() // U+3FC9 <cjk>
	0x88: [`\u7641`].string() // U+7641 <cjk>
	0x89: utf32_to_str(0x24E8B) // U+24E8B <cjk>
	0x8A: [`\u7649`].string() // U+7649 <cjk>
	0x8B: [`\u7655`].string() // U+7655 <cjk>
	0x8C: [`\u3FD7`].string() // U+3FD7 <cjk>
	0x8D: [`\u766E`].string() // U+766E <cjk>
	0x8E: [`\u7695`].string() // U+7695 <cjk>
	0x8F: [`\u769C`].string() // U+769C <cjk>
	0x90: [`\u76A1`].string() // U+76A1 <cjk>
	0x91: [`\u76A0`].string() // U+76A0 <cjk>
	0x92: [`\u76A7`].string() // U+76A7 <cjk>
	0x93: [`\u76A8`].string() // U+76A8 <cjk>
	0x94: [`\u76AF`].string() // U+76AF <cjk>
	0x95: utf32_to_str(0x2504A) // U+2504A <cjk>
	0x96: [`\u76C9`].string() // U+76C9 <cjk>
	0x97: utf32_to_str(0x25055) // U+25055 <cjk>
	0x98: [`\u76E8`].string() // U+76E8 <cjk>
	0x99: [`\u76EC`].string() // U+76EC <cjk>
	0x9A: utf32_to_str(0x25122) // U+25122 <cjk>
	0x9B: [`\u7717`].string() // U+7717 <cjk>
	0x9C: [`\u771A`].string() // U+771A <cjk>
	0x9D: [`\u772D`].string() // U+772D <cjk>
	0x9E: [`\u7735`].string() // U+7735 <cjk>
	0x9F: utf32_to_str(0x251A9) // U+251A9 <cjk>
	0xA0: [`\u4039`].string() // U+4039 <cjk>
	0xA1: utf32_to_str(0x251E5) // U+251E5 <cjk>
	0xA2: utf32_to_str(0x251CD) // U+251CD <cjk>
	0xA3: [`\u7758`].string() // U+7758 <cjk>
	0xA4: [`\u7760`].string() // U+7760 <cjk>
	0xA5: [`\u776A`].string() // U+776A <cjk>
	0xA6: utf32_to_str(0x2521E) // U+2521E <cjk>
	0xA7: [`\u7772`].string() // U+7772 <cjk>
	0xA8: [`\u777C`].string() // U+777C <cjk>
	0xA9: [`\u777D`].string() // U+777D <cjk>
	0xAA: utf32_to_str(0x2524C) // U+2524C <cjk>
	0xAB: [`\u4058`].string() // U+4058 <cjk>
	0xAC: [`\u779A`].string() // U+779A <cjk>
	0xAD: [`\u779F`].string() // U+779F <cjk>
	0xAE: [`\u77A2`].string() // U+77A2 <cjk>
	0xAF: [`\u77A4`].string() // U+77A4 <cjk>
	0xB0: [`\u77A9`].string() // U+77A9 <cjk>
	0xB1: [`\u77DE`].string() // U+77DE <cjk>
	0xB2: [`\u77DF`].string() // U+77DF <cjk>
	0xB3: [`\u77E4`].string() // U+77E4 <cjk>
	0xB4: [`\u77E6`].string() // U+77E6 <cjk>
	0xB5: [`\u77EA`].string() // U+77EA <cjk>
	0xB6: [`\u77EC`].string() // U+77EC <cjk>
	0xB7: [`\u4093`].string() // U+4093 <cjk>
	0xB8: [`\u77F0`].string() // U+77F0 <cjk>
	0xB9: [`\u77F4`].string() // U+77F4 <cjk>
	0xBA: [`\u77FB`].string() // U+77FB <cjk>
	0xBB: utf32_to_str(0x2542E) // U+2542E <cjk>
	0xBC: [`\u7805`].string() // U+7805 <cjk>
	0xBD: [`\u7806`].string() // U+7806 <cjk>
	0xBE: [`\u7809`].string() // U+7809 <cjk>
	0xBF: [`\u780D`].string() // U+780D <cjk>
	0xC0: [`\u7819`].string() // U+7819 <cjk>
	0xC1: [`\u7821`].string() // U+7821 <cjk>
	0xC2: [`\u782C`].string() // U+782C <cjk>
	0xC3: [`\u7847`].string() // U+7847 <cjk>
	0xC4: [`\u7864`].string() // U+7864 <cjk>
	0xC5: [`\u786A`].string() // U+786A <cjk>
	0xC6: utf32_to_str(0x254D9) // U+254D9 <cjk>
	0xC7: [`\u788A`].string() // U+788A <cjk>
	0xC8: [`\u7894`].string() // U+7894 <cjk>
	0xC9: [`\u78A4`].string() // U+78A4 <cjk>
	0xCA: [`\u789D`].string() // U+789D <cjk>
	0xCB: [`\u789E`].string() // U+789E <cjk>
	0xCC: [`\u789F`].string() // U+789F <cjk>
	0xCD: [`\u78BB`].string() // U+78BB <cjk>
	0xCE: [`\u78C8`].string() // U+78C8 <cjk>
	0xCF: [`\u78CC`].string() // U+78CC <cjk>
	0xD0: [`\u78CE`].string() // U+78CE <cjk>
	0xD1: [`\u78D5`].string() // U+78D5 <cjk>
	0xD2: [`\u78E0`].string() // U+78E0 <cjk>
	0xD3: [`\u78E1`].string() // U+78E1 <cjk>
	0xD4: [`\u78E6`].string() // U+78E6 <cjk>
	0xD5: [`\u78F9`].string() // U+78F9 <cjk>
	0xD6: [`\u78FA`].string() // U+78FA <cjk>
	0xD7: [`\u78FB`].string() // U+78FB <cjk>
	0xD8: [`\u78FE`].string() // U+78FE <cjk>
	0xD9: utf32_to_str(0x255A7) // U+255A7 <cjk>
	0xDA: [`\u7910`].string() // U+7910 <cjk>
	0xDB: [`\u791B`].string() // U+791B <cjk>
	0xDC: [`\u7930`].string() // U+7930 <cjk>
	0xDD: [`\u7925`].string() // U+7925 <cjk>
	0xDE: [`\u793B`].string() // U+793B <cjk>
	0xDF: [`\u794A`].string() // U+794A <cjk>
	0xE0: [`\u7958`].string() // U+7958 <cjk>
	0xE1: [`\u795B`].string() // U+795B <cjk>
	0xE2: [`\u4105`].string() // U+4105 <cjk>
	0xE3: [`\u7967`].string() // U+7967 <cjk>
	0xE4: [`\u7972`].string() // U+7972 <cjk>
	0xE5: [`\u7994`].string() // U+7994 <cjk>
	0xE6: [`\u7995`].string() // U+7995 <cjk>
	0xE7: [`\u7996`].string() // U+7996 <cjk>
	0xE8: [`\u799B`].string() // U+799B <cjk>
	0xE9: [`\u79A1`].string() // U+79A1 <cjk>
	0xEA: [`\u79A9`].string() // U+79A9 <cjk>
	0xEB: [`\u79B4`].string() // U+79B4 <cjk>
	0xEC: [`\u79BB`].string() // U+79BB <cjk>
	0xED: [`\u79C2`].string() // U+79C2 <cjk>
	0xEE: [`\u79C7`].string() // U+79C7 <cjk>
	0xEF: [`\u79CC`].string() // U+79CC <cjk>
	0xF0: [`\u79CD`].string() // U+79CD <cjk>
	0xF1: [`\u79D6`].string() // U+79D6 <cjk>
	0xF2: [`\u4148`].string() // U+4148 <cjk>
	0xF3: utf32_to_str(0x257A9) // U+257A9 <cjk>
	0xF4: utf32_to_str(0x257B4) // U+257B4 <cjk>
	0xF5: [`\u414F`].string() // U+414F <cjk>
	0xF6: [`\u7A0A`].string() // U+7A0A <cjk>
	0xF7: [`\u7A11`].string() // U+7A11 <cjk>
	0xF8: [`\u7A15`].string() // U+7A15 <cjk>
	0xF9: [`\u7A1B`].string() // U+7A1B <cjk>
	0xFA: [`\u7A1E`].string() // U+7A1E <cjk>
	0xFB: [`\u4163`].string() // U+4163 <cjk>
	0xFC: [`\u7A2D`].string() // U+7A2D <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xf1 = {
	0x40: [`\u5108`].string() // U+5108 <cjk>
	0x41: utf32_to_str(0x203F9) // U+203F9 <cjk>
	0x42: [`\u5117`].string() // U+5117 <cjk>
	0x43: [`\u511B`].string() // U+511B <cjk>
	0x44: utf32_to_str(0x2044A) // U+2044A <cjk>
	0x45: [`\u5160`].string() // U+5160 <cjk>
	0x46: utf32_to_str(0x20509) // U+20509 <cjk>
	0x47: [`\u5173`].string() // U+5173 <cjk>
	0x48: [`\u5183`].string() // U+5183 <cjk>
	0x49: [`\u518B`].string() // U+518B <cjk>
	0x4A: [`\u34BC`].string() // U+34BC <cjk>
	0x4B: [`\u5198`].string() // U+5198 <cjk>
	0x4C: [`\u51A3`].string() // U+51A3 <cjk>
	0x4D: [`\u51AD`].string() // U+51AD <cjk>
	0x4E: [`\u34C7`].string() // U+34C7 <cjk>
	0x4F: [`\u51BC`].string() // U+51BC <cjk>
	0x50: utf32_to_str(0x205D6) // U+205D6 <cjk>
	0x51: utf32_to_str(0x20628) // U+20628 <cjk>
	0x52: [`\u51F3`].string() // U+51F3 <cjk>
	0x53: [`\u51F4`].string() // U+51F4 <cjk>
	0x54: [`\u5202`].string() // U+5202 <cjk>
	0x55: [`\u5212`].string() // U+5212 <cjk>
	0x56: [`\u5216`].string() // U+5216 <cjk>
	0x57: utf32_to_str(0x2074F) // U+2074F <cjk>
	0x58: [`\u5255`].string() // U+5255 <cjk>
	0x59: [`\u525C`].string() // U+525C <cjk>
	0x5A: [`\u526C`].string() // U+526C <cjk>
	0x5B: [`\u5277`].string() // U+5277 <cjk>
	0x5C: [`\u5284`].string() // U+5284 <cjk>
	0x5D: [`\u5282`].string() // U+5282 <cjk>
	0x5E: utf32_to_str(0x20807) // U+20807 <cjk>
	0x5F: [`\u5298`].string() // U+5298 <cjk>
	0x60: utf32_to_str(0x2083A) // U+2083A <cjk>
	0x61: [`\u52A4`].string() // U+52A4 <cjk>
	0x62: [`\u52A6`].string() // U+52A6 <cjk>
	0x63: [`\u52AF`].string() // U+52AF <cjk>
	0x64: [`\u52BA`].string() // U+52BA <cjk>
	0x65: [`\u52BB`].string() // U+52BB <cjk>
	0x66: [`\u52CA`].string() // U+52CA <cjk>
	0x67: [`\u351F`].string() // U+351F <cjk>
	0x68: [`\u52D1`].string() // U+52D1 <cjk>
	0x69: utf32_to_str(0x208B9) // U+208B9 <cjk>
	0x6A: [`\u52F7`].string() // U+52F7 <cjk>
	0x6B: [`\u530A`].string() // U+530A <cjk>
	0x6C: [`\u530B`].string() // U+530B <cjk>
	0x6D: [`\u5324`].string() // U+5324 <cjk>
	0x6E: [`\u5335`].string() // U+5335 <cjk>
	0x6F: [`\u533E`].string() // U+533E <cjk>
	0x70: [`\u5342`].string() // U+5342 <cjk>
	0x71: utf32_to_str(0x2097C) // U+2097C <cjk>
	0x72: utf32_to_str(0x2099D) // U+2099D <cjk>
	0x73: [`\u5367`].string() // U+5367 <cjk>
	0x74: [`\u536C`].string() // U+536C <cjk>
	0x75: [`\u537A`].string() // U+537A <cjk>
	0x76: [`\u53A4`].string() // U+53A4 <cjk>
	0x77: [`\u53B4`].string() // U+53B4 <cjk>
	0x78: utf32_to_str(0x20AD3) // U+20AD3 <cjk>
	0x79: [`\u53B7`].string() // U+53B7 <cjk>
	0x7A: [`\u53C0`].string() // U+53C0 <cjk>
	0x7B: utf32_to_str(0x20B1D) // U+20B1D <cjk>
	0x7C: [`\u355D`].string() // U+355D <cjk>
	0x7D: [`\u355E`].string() // U+355E <cjk>
	0x7E: [`\u53D5`].string() // U+53D5 <cjk>
	0x80: [`\u53DA`].string() // U+53DA <cjk>
	0x81: [`\u3563`].string() // U+3563 <cjk>
	0x82: [`\u53F4`].string() // U+53F4 <cjk>
	0x83: [`\u53F5`].string() // U+53F5 <cjk>
	0x84: [`\u5455`].string() // U+5455 <cjk>
	0x85: [`\u5424`].string() // U+5424 <cjk>
	0x86: [`\u5428`].string() // U+5428 <cjk>
	0x87: [`\u356E`].string() // U+356E <cjk>
	0x88: [`\u5443`].string() // U+5443 <cjk>
	0x89: [`\u5462`].string() // U+5462 <cjk>
	0x8A: [`\u5466`].string() // U+5466 <cjk>
	0x8B: [`\u546C`].string() // U+546C <cjk>
	0x8C: [`\u548A`].string() // U+548A <cjk>
	0x8D: [`\u548D`].string() // U+548D <cjk>
	0x8E: [`\u5495`].string() // U+5495 <cjk>
	0x8F: [`\u54A0`].string() // U+54A0 <cjk>
	0x90: [`\u54A6`].string() // U+54A6 <cjk>
	0x91: [`\u54AD`].string() // U+54AD <cjk>
	0x92: [`\u54AE`].string() // U+54AE <cjk>
	0x93: [`\u54B7`].string() // U+54B7 <cjk>
	0x94: [`\u54BA`].string() // U+54BA <cjk>
	0x95: [`\u54BF`].string() // U+54BF <cjk>
	0x96: [`\u54C3`].string() // U+54C3 <cjk>
	0x97: utf32_to_str(0x20D45) // U+20D45 <cjk>
	0x98: [`\u54EC`].string() // U+54EC <cjk>
	0x99: [`\u54EF`].string() // U+54EF <cjk>
	0x9A: [`\u54F1`].string() // U+54F1 <cjk>
	0x9B: [`\u54F3`].string() // U+54F3 <cjk>
	0x9C: [`\u5500`].string() // U+5500 <cjk>
	0x9D: [`\u5501`].string() // U+5501 <cjk>
	0x9E: [`\u5509`].string() // U+5509 <cjk>
	0x9F: [`\u553C`].string() // U+553C <cjk>
	0xA0: [`\u5541`].string() // U+5541 <cjk>
	0xA1: [`\u35A6`].string() // U+35A6 <cjk>
	0xA2: [`\u5547`].string() // U+5547 <cjk>
	0xA3: [`\u554A`].string() // U+554A <cjk>
	0xA4: [`\u35A8`].string() // U+35A8 <cjk>
	0xA5: [`\u5560`].string() // U+5560 <cjk>
	0xA6: [`\u5561`].string() // U+5561 <cjk>
	0xA7: [`\u5564`].string() // U+5564 <cjk>
	0xA8: utf32_to_str(0x20DE1) // U+20DE1 <cjk>
	0xA9: [`\u557D`].string() // U+557D <cjk>
	0xAA: [`\u5582`].string() // U+5582 <cjk>
	0xAB: [`\u5588`].string() // U+5588 <cjk>
	0xAC: [`\u5591`].string() // U+5591 <cjk>
	0xAD: [`\u35C5`].string() // U+35C5 <cjk>
	0xAE: [`\u55D2`].string() // U+55D2 <cjk>
	0xAF: utf32_to_str(0x20E95) // U+20E95 <cjk>
	0xB0: utf32_to_str(0x20E6D) // U+20E6D <cjk>
	0xB1: [`\u55BF`].string() // U+55BF <cjk>
	0xB2: [`\u55C9`].string() // U+55C9 <cjk>
	0xB3: [`\u55CC`].string() // U+55CC <cjk>
	0xB4: [`\u55D1`].string() // U+55D1 <cjk>
	0xB5: [`\u55DD`].string() // U+55DD <cjk>
	0xB6: [`\u35DA`].string() // U+35DA <cjk>
	0xB7: [`\u55E2`].string() // U+55E2 <cjk>
	0xB8: utf32_to_str(0x20E64) // U+20E64 <cjk>
	0xB9: [`\u55E9`].string() // U+55E9 <cjk>
	0xBA: [`\u5628`].string() // U+5628 <cjk>
	0xBB: utf32_to_str(0x20F5F) // U+20F5F <cjk>
	0xBC: [`\u5607`].string() // U+5607 <cjk>
	0xBD: [`\u5610`].string() // U+5610 <cjk>
	0xBE: [`\u5630`].string() // U+5630 <cjk>
	0xBF: [`\u5637`].string() // U+5637 <cjk>
	0xC0: [`\u35F4`].string() // U+35F4 <cjk>
	0xC1: [`\u563D`].string() // U+563D <cjk>
	0xC2: [`\u563F`].string() // U+563F <cjk>
	0xC3: [`\u5640`].string() // U+5640 <cjk>
	0xC4: [`\u5647`].string() // U+5647 <cjk>
	0xC5: [`\u565E`].string() // U+565E <cjk>
	0xC6: [`\u5660`].string() // U+5660 <cjk>
	0xC7: [`\u566D`].string() // U+566D <cjk>
	0xC8: [`\u3605`].string() // U+3605 <cjk>
	0xC9: [`\u5688`].string() // U+5688 <cjk>
	0xCA: [`\u568C`].string() // U+568C <cjk>
	0xCB: [`\u5695`].string() // U+5695 <cjk>
	0xCC: [`\u569A`].string() // U+569A <cjk>
	0xCD: [`\u569D`].string() // U+569D <cjk>
	0xCE: [`\u56A8`].string() // U+56A8 <cjk>
	0xCF: [`\u56AD`].string() // U+56AD <cjk>
	0xD0: [`\u56B2`].string() // U+56B2 <cjk>
	0xD1: [`\u56C5`].string() // U+56C5 <cjk>
	0xD2: [`\u56CD`].string() // U+56CD <cjk>
	0xD3: [`\u56DF`].string() // U+56DF <cjk>
	0xD4: [`\u56E8`].string() // U+56E8 <cjk>
	0xD5: [`\u56F6`].string() // U+56F6 <cjk>
	0xD6: [`\u56F7`].string() // U+56F7 <cjk>
	0xD7: utf32_to_str(0x21201) // U+21201 <cjk>
	0xD8: [`\u5715`].string() // U+5715 <cjk>
	0xD9: [`\u5723`].string() // U+5723 <cjk>
	0xDA: utf32_to_str(0x21255) // U+21255 <cjk>
	0xDB: [`\u5729`].string() // U+5729 <cjk>
	0xDC: utf32_to_str(0x2127B) // U+2127B <cjk>
	0xDD: [`\u5745`].string() // U+5745 <cjk>
	0xDE: [`\u5746`].string() // U+5746 <cjk>
	0xDF: [`\u574C`].string() // U+574C <cjk>
	0xE0: [`\u574D`].string() // U+574D <cjk>
	0xE1: utf32_to_str(0x21274) // U+21274 <cjk>
	0xE2: [`\u5768`].string() // U+5768 <cjk>
	0xE3: [`\u576F`].string() // U+576F <cjk>
	0xE4: [`\u5773`].string() // U+5773 <cjk>
	0xE5: [`\u5774`].string() // U+5774 <cjk>
	0xE6: [`\u5775`].string() // U+5775 <cjk>
	0xE7: [`\u577B`].string() // U+577B <cjk>
	0xE8: utf32_to_str(0x212E4) // U+212E4 <cjk>
	0xE9: utf32_to_str(0x212D7) // U+212D7 <cjk>
	0xEA: [`\u57AC`].string() // U+57AC <cjk>
	0xEB: [`\u579A`].string() // U+579A <cjk>
	0xEC: [`\u579D`].string() // U+579D <cjk>
	0xED: [`\u579E`].string() // U+579E <cjk>
	0xEE: [`\u57A8`].string() // U+57A8 <cjk>
	0xEF: [`\u57D7`].string() // U+57D7 <cjk>
	0xF0: utf32_to_str(0x212FD) // U+212FD <cjk>
	0xF1: [`\u57CC`].string() // U+57CC <cjk>
	0xF2: utf32_to_str(0x21336) // U+21336 <cjk>
	0xF3: utf32_to_str(0x21344) // U+21344 <cjk>
	0xF4: [`\u57DE`].string() // U+57DE <cjk>
	0xF5: [`\u57E6`].string() // U+57E6 <cjk>
	0xF6: [`\u57F0`].string() // U+57F0 <cjk>
	0xF7: [`\u364A`].string() // U+364A <cjk>
	0xF8: [`\u57F8`].string() // U+57F8 <cjk>
	0xF9: [`\u57FB`].string() // U+57FB <cjk>
	0xFA: [`\u57FD`].string() // U+57FD <cjk>
	0xFB: [`\u5804`].string() // U+5804 <cjk>
	0xFC: [`\u581E`].string() // U+581E <cjk>
}

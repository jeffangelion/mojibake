module mojibake

const jis_x_0213_doublebyte_0x99 = {
	0x40: [`\u50C9`].string() // U+50C9 <cjk>
	0x41: [`\u50CA`].string() // U+50CA <cjk>
	0x42: [`\u50B3`].string() // U+50B3 <cjk>
	0x43: [`\u50C2`].string() // U+50C2 <cjk>
	0x44: [`\u50D6`].string() // U+50D6 <cjk>
	0x45: [`\u50DE`].string() // U+50DE <cjk>
	0x46: [`\u50E5`].string() // U+50E5 <cjk>
	0x47: [`\u50ED`].string() // U+50ED <cjk>
	0x48: [`\u50E3`].string() // U+50E3 <cjk>
	0x49: [`\u50EE`].string() // U+50EE <cjk>
	0x4A: [`\u50F9`].string() // U+50F9 <cjk>
	0x4B: [`\u50F5`].string() // U+50F5 <cjk>
	0x4C: [`\u5109`].string() // U+5109 <cjk>
	0x4D: [`\u5101`].string() // U+5101 <cjk>
	0x4E: [`\u5102`].string() // U+5102 <cjk>
	0x4F: [`\u5116`].string() // U+5116 <cjk>
	0x50: [`\u5115`].string() // U+5115 <cjk>
	0x51: [`\u5114`].string() // U+5114 <cjk>
	0x52: [`\u511A`].string() // U+511A <cjk>
	0x53: [`\u5121`].string() // U+5121 <cjk>
	0x54: [`\u513A`].string() // U+513A <cjk>
	0x55: [`\u5137`].string() // U+5137 <cjk>
	0x56: [`\u513C`].string() // U+513C <cjk>
	0x57: [`\u513B`].string() // U+513B <cjk>
	0x58: [`\u513F`].string() // U+513F <cjk>
	0x59: [`\u5140`].string() // U+5140 <cjk>
	0x5A: [`\u5152`].string() // U+5152 <cjk>
	0x5B: [`\u514C`].string() // U+514C <cjk>
	0x5C: [`\u5154`].string() // U+5154 <cjk>
	0x5D: [`\u5162`].string() // U+5162 <cjk>
	0x5E: [`\u7AF8`].string() // U+7AF8 <cjk>
	0x5F: [`\u5169`].string() // U+5169 <cjk>
	0x60: [`\u516A`].string() // U+516A <cjk>
	0x61: [`\u516E`].string() // U+516E <cjk>
	0x62: [`\u5180`].string() // U+5180 <cjk>
	0x63: [`\u5182`].string() // U+5182 <cjk>
	0x64: [`\u56D8`].string() // U+56D8 <cjk>
	0x65: [`\u518C`].string() // U+518C <cjk>
	0x66: [`\u5189`].string() // U+5189 <cjk>
	0x67: [`\u518F`].string() // U+518F <cjk>
	0x68: [`\u5191`].string() // U+5191 <cjk>
	0x69: [`\u5193`].string() // U+5193 <cjk>
	0x6A: [`\u5195`].string() // U+5195 <cjk>
	0x6B: [`\u5196`].string() // U+5196 <cjk>
	0x6C: [`\u51A4`].string() // U+51A4 <cjk>
	0x6D: [`\u51A6`].string() // U+51A6 <cjk>
	0x6E: [`\u51A2`].string() // U+51A2 <cjk>
	0x6F: [`\u51A9`].string() // U+51A9 <cjk>
	0x70: [`\u51AA`].string() // U+51AA <cjk>
	0x71: [`\u51AB`].string() // U+51AB <cjk>
	0x72: [`\u51B3`].string() // U+51B3 <cjk>
	0x73: [`\u51B1`].string() // U+51B1 <cjk>
	0x74: [`\u51B2`].string() // U+51B2 <cjk>
	0x75: [`\u51B0`].string() // U+51B0 <cjk>
	0x76: [`\u51B5`].string() // U+51B5 <cjk>
	0x77: [`\u51BD`].string() // U+51BD <cjk>
	0x78: [`\u51C5`].string() // U+51C5 <cjk>
	0x79: [`\u51C9`].string() // U+51C9 <cjk>
	0x7A: [`\u51DB`].string() // U+51DB <cjk>
	0x7B: [`\u51E0`].string() // U+51E0 <cjk>
	0x7C: [`\u8655`].string() // U+8655 <cjk>
	0x7D: [`\u51E9`].string() // U+51E9 <cjk>
	0x7E: [`\u51ED`].string() // U+51ED <cjk>
	0x80: [`\u51F0`].string() // U+51F0 <cjk>
	0x81: [`\u51F5`].string() // U+51F5 <cjk>
	0x82: [`\u51FE`].string() // U+51FE <cjk>
	0x83: [`\u5204`].string() // U+5204 <cjk>
	0x84: [`\u520B`].string() // U+520B <cjk>
	0x85: [`\u5214`].string() // U+5214 <cjk>
	0x86: [`\u520E`].string() // U+520E <cjk>
	0x87: [`\u5227`].string() // U+5227 <cjk>
	0x88: [`\u522A`].string() // U+522A <cjk>
	0x89: [`\u522E`].string() // U+522E <cjk>
	0x8A: [`\u5233`].string() // U+5233 <cjk>
	0x8B: [`\u5239`].string() // U+5239 <cjk>
	0x8C: [`\u524F`].string() // U+524F <cjk>
	0x8D: [`\u5244`].string() // U+5244 <cjk>
	0x8E: [`\u524B`].string() // U+524B <cjk>
	0x8F: [`\u524C`].string() // U+524C <cjk>
	0x90: [`\u525E`].string() // U+525E <cjk>
	0x91: [`\u5254`].string() // U+5254 <cjk>
	0x92: [`\u526A`].string() // U+526A <cjk>
	0x93: [`\u5274`].string() // U+5274 <cjk>
	0x94: [`\u5269`].string() // U+5269 <cjk>
	0x95: [`\u5273`].string() // U+5273 <cjk>
	0x96: [`\u527F`].string() // U+527F <cjk>
	0x97: [`\u527D`].string() // U+527D <cjk>
	0x98: [`\u528D`].string() // U+528D <cjk>
	0x99: [`\u5294`].string() // U+5294 <cjk>
	0x9A: [`\u5292`].string() // U+5292 <cjk>
	0x9B: [`\u5271`].string() // U+5271 <cjk>
	0x9C: [`\u5288`].string() // U+5288 <cjk>
	0x9D: [`\u5291`].string() // U+5291 <cjk>
	0x9E: [`\u8FA8`].string() // U+8FA8 <cjk>
	0x9F: [`\u8FA7`].string() // U+8FA7 <cjk>
	0xA0: [`\u52AC`].string() // U+52AC <cjk>
	0xA1: [`\u52AD`].string() // U+52AD <cjk>
	0xA2: [`\u52BC`].string() // U+52BC <cjk>
	0xA3: [`\u52B5`].string() // U+52B5 <cjk>
	0xA4: [`\u52C1`].string() // U+52C1 <cjk>
	0xA5: [`\u52CD`].string() // U+52CD <cjk>
	0xA6: [`\u52D7`].string() // U+52D7 <cjk>
	0xA7: [`\u52DE`].string() // U+52DE <cjk>
	0xA8: [`\u52E3`].string() // U+52E3 <cjk>
	0xA9: [`\u52E6`].string() // U+52E6 <cjk>
	0xAA: [`\u98ED`].string() // U+98ED <cjk>
	0xAB: [`\u52E0`].string() // U+52E0 <cjk>
	0xAC: [`\u52F3`].string() // U+52F3 <cjk>
	0xAD: [`\u52F5`].string() // U+52F5 <cjk>
	0xAE: [`\u52F8`].string() // U+52F8 <cjk>
	0xAF: [`\u52F9`].string() // U+52F9 <cjk>
	0xB0: [`\u5306`].string() // U+5306 <cjk>
	0xB1: [`\u5308`].string() // U+5308 <cjk>
	0xB2: [`\u7538`].string() // U+7538 <cjk>
	0xB3: [`\u530D`].string() // U+530D <cjk>
	0xB4: [`\u5310`].string() // U+5310 <cjk>
	0xB5: [`\u530F`].string() // U+530F <cjk>
	0xB6: [`\u5315`].string() // U+5315 <cjk>
	0xB7: [`\u531A`].string() // U+531A <cjk>
	0xB8: [`\u5323`].string() // U+5323 <cjk>
	0xB9: [`\u532F`].string() // U+532F <cjk>
	0xBA: [`\u5331`].string() // U+5331 <cjk>
	0xBB: [`\u5333`].string() // U+5333 <cjk>
	0xBC: [`\u5338`].string() // U+5338 <cjk>
	0xBD: [`\u5340`].string() // U+5340 <cjk>
	0xBE: [`\u5346`].string() // U+5346 <cjk>
	0xBF: [`\u5345`].string() // U+5345 <cjk>
	0xC0: [`\u4E17`].string() // U+4E17 <cjk>
	0xC1: [`\u5349`].string() // U+5349 <cjk>
	0xC2: [`\u534D`].string() // U+534D <cjk>
	0xC3: [`\u51D6`].string() // U+51D6 <cjk>
	0xC4: [`\u535E`].string() // U+535E <cjk>
	0xC5: [`\u5369`].string() // U+5369 <cjk>
	0xC6: [`\u536E`].string() // U+536E <cjk>
	0xC7: [`\u5918`].string() // U+5918 <cjk>
	0xC8: [`\u537B`].string() // U+537B <cjk>
	0xC9: [`\u5377`].string() // U+5377 <cjk>
	0xCA: [`\u5382`].string() // U+5382 <cjk>
	0xCB: [`\u5396`].string() // U+5396 <cjk>
	0xCC: [`\u53A0`].string() // U+53A0 <cjk>
	0xCD: [`\u53A6`].string() // U+53A6 <cjk>
	0xCE: [`\u53A5`].string() // U+53A5 <cjk>
	0xCF: [`\u53AE`].string() // U+53AE <cjk>
	0xD0: [`\u53B0`].string() // U+53B0 <cjk>
	0xD1: [`\u53B6`].string() // U+53B6 <cjk>
	0xD2: [`\u53C3`].string() // U+53C3 <cjk>
	0xD3: [`\u7C12`].string() // U+7C12 <cjk>
	0xD4: [`\u96D9`].string() // U+96D9 <cjk>
	0xD5: [`\u53DF`].string() // U+53DF <cjk>
	0xD6: [`\u66FC`].string() // U+66FC <cjk>
	0xD7: [`\u71EE`].string() // U+71EE <cjk>
	0xD8: [`\u53EE`].string() // U+53EE <cjk>
	0xD9: [`\u53E8`].string() // U+53E8 <cjk>
	0xDA: [`\u53ED`].string() // U+53ED <cjk>
	0xDB: [`\u53FA`].string() // U+53FA <cjk>
	0xDC: [`\u5401`].string() // U+5401 <cjk>
	0xDD: [`\u543D`].string() // U+543D <cjk>
	0xDE: [`\u5440`].string() // U+5440 <cjk>
	0xDF: [`\u542C`].string() // U+542C <cjk>
	0xE0: [`\u542D`].string() // U+542D <cjk>
	0xE1: [`\u543C`].string() // U+543C <cjk>
	0xE2: [`\u542E`].string() // U+542E <cjk>
	0xE3: [`\u5436`].string() // U+5436 <cjk>
	0xE4: [`\u5429`].string() // U+5429 <cjk>
	0xE5: [`\u541D`].string() // U+541D <cjk>
	0xE6: [`\u544E`].string() // U+544E <cjk>
	0xE7: [`\u548F`].string() // U+548F <cjk>
	0xE8: [`\u5475`].string() // U+5475 <cjk>
	0xE9: [`\u548E`].string() // U+548E <cjk>
	0xEA: [`\u545F`].string() // U+545F <cjk>
	0xEB: [`\u5471`].string() // U+5471 <cjk>
	0xEC: [`\u5477`].string() // U+5477 <cjk>
	0xED: [`\u5470`].string() // U+5470 <cjk>
	0xEE: [`\u5492`].string() // U+5492 <cjk>
	0xEF: [`\u547B`].string() // U+547B <cjk>
	0xF0: [`\u5480`].string() // U+5480 <cjk>
	0xF1: [`\u5476`].string() // U+5476 <cjk>
	0xF2: [`\u5484`].string() // U+5484 <cjk>
	0xF3: [`\u5490`].string() // U+5490 <cjk>
	0xF4: [`\u5486`].string() // U+5486 <cjk>
	0xF5: [`\u54C7`].string() // U+54C7 <cjk>
	0xF6: [`\u54A2`].string() // U+54A2 <cjk>
	0xF7: [`\u54B8`].string() // U+54B8 <cjk>
	0xF8: [`\u54A5`].string() // U+54A5 <cjk>
	0xF9: [`\u54AC`].string() // U+54AC <cjk>
	0xFA: [`\u54C4`].string() // U+54C4 <cjk>
	0xFB: [`\u54C8`].string() // U+54C8 <cjk>
	0xFC: [`\u54A8`].string() // U+54A8 <cjk>
}

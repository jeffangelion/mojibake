module mojibake

const jis_x_0213_doublebyte_0xf5 = {
	0x40: [`\u6E93`].string() // U+6E93 <cjk>
	0x41: [`\u6EA7`].string() // U+6EA7 <cjk>
	0x42: [`\u6EB4`].string() // U+6EB4 <cjk>
	0x43: [`\u6EBF`].string() // U+6EBF <cjk>
	0x44: [`\u6EC3`].string() // U+6EC3 <cjk>
	0x45: [`\u6ECA`].string() // U+6ECA <cjk>
	0x46: [`\u6ED9`].string() // U+6ED9 <cjk>
	0x47: [`\u6F35`].string() // U+6F35 <cjk>
	0x48: [`\u6EEB`].string() // U+6EEB <cjk>
	0x49: [`\u6EF9`].string() // U+6EF9 <cjk>
	0x4A: [`\u6EFB`].string() // U+6EFB <cjk>
	0x4B: [`\u6F0A`].string() // U+6F0A <cjk>
	0x4C: [`\u6F0C`].string() // U+6F0C <cjk>
	0x4D: [`\u6F18`].string() // U+6F18 <cjk>
	0x4E: [`\u6F25`].string() // U+6F25 <cjk>
	0x4F: [`\u6F36`].string() // U+6F36 <cjk>
	0x50: [`\u6F3C`].string() // U+6F3C <cjk>
	0x51: utf32_to_str(0x23F7E) // U+23F7E <cjk>
	0x52: [`\u6F52`].string() // U+6F52 <cjk>
	0x53: [`\u6F57`].string() // U+6F57 <cjk>
	0x54: [`\u6F5A`].string() // U+6F5A <cjk>
	0x55: [`\u6F60`].string() // U+6F60 <cjk>
	0x56: [`\u6F68`].string() // U+6F68 <cjk>
	0x57: [`\u6F98`].string() // U+6F98 <cjk>
	0x58: [`\u6F7D`].string() // U+6F7D <cjk>
	0x59: [`\u6F90`].string() // U+6F90 <cjk>
	0x5A: [`\u6F96`].string() // U+6F96 <cjk>
	0x5B: [`\u6FBE`].string() // U+6FBE <cjk>
	0x5C: [`\u6F9F`].string() // U+6F9F <cjk>
	0x5D: [`\u6FA5`].string() // U+6FA5 <cjk>
	0x5E: [`\u6FAF`].string() // U+6FAF <cjk>
	0x5F: [`\u3D64`].string() // U+3D64 <cjk>
	0x60: [`\u6FB5`].string() // U+6FB5 <cjk>
	0x61: [`\u6FC8`].string() // U+6FC8 <cjk>
	0x62: [`\u6FC9`].string() // U+6FC9 <cjk>
	0x63: [`\u6FDA`].string() // U+6FDA <cjk>
	0x64: [`\u6FDE`].string() // U+6FDE <cjk>
	0x65: [`\u6FE9`].string() // U+6FE9 <cjk>
	0x66: utf32_to_str(0x24096) // U+24096 <cjk>
	0x67: [`\u6FFC`].string() // U+6FFC <cjk>
	0x68: [`\u7000`].string() // U+7000 <cjk>
	0x69: [`\u7007`].string() // U+7007 <cjk>
	0x6A: [`\u700A`].string() // U+700A <cjk>
	0x6B: [`\u7023`].string() // U+7023 <cjk>
	0x6C: utf32_to_str(0x24103) // U+24103 <cjk>
	0x6D: [`\u7039`].string() // U+7039 <cjk>
	0x6E: [`\u703A`].string() // U+703A <cjk>
	0x6F: [`\u703C`].string() // U+703C <cjk>
	0x70: [`\u7043`].string() // U+7043 <cjk>
	0x71: [`\u7047`].string() // U+7047 <cjk>
	0x72: [`\u704B`].string() // U+704B <cjk>
	0x73: [`\u3D9A`].string() // U+3D9A <cjk>
	0x74: [`\u7054`].string() // U+7054 <cjk>
	0x75: [`\u7065`].string() // U+7065 <cjk>
	0x76: [`\u7069`].string() // U+7069 <cjk>
	0x77: [`\u706C`].string() // U+706C <cjk>
	0x78: [`\u706E`].string() // U+706E <cjk>
	0x79: [`\u7076`].string() // U+7076 <cjk>
	0x7A: [`\u707E`].string() // U+707E <cjk>
	0x7B: [`\u7081`].string() // U+7081 <cjk>
	0x7C: [`\u7086`].string() // U+7086 <cjk>
	0x7D: [`\u7095`].string() // U+7095 <cjk>
	0x7E: [`\u7097`].string() // U+7097 <cjk>
	0x80: [`\u70BB`].string() // U+70BB <cjk>
	0x81: utf32_to_str(0x241C6) // U+241C6 <cjk>
	0x82: [`\u709F`].string() // U+709F <cjk>
	0x83: [`\u70B1`].string() // U+70B1 <cjk>
	0x84: utf32_to_str(0x241FE) // U+241FE <cjk>
	0x85: [`\u70EC`].string() // U+70EC <cjk>
	0x86: [`\u70CA`].string() // U+70CA <cjk>
	0x87: [`\u70D1`].string() // U+70D1 <cjk>
	0x88: [`\u70D3`].string() // U+70D3 <cjk>
	0x89: [`\u70DC`].string() // U+70DC <cjk>
	0x8A: [`\u7103`].string() // U+7103 <cjk>
	0x8B: [`\u7104`].string() // U+7104 <cjk>
	0x8C: [`\u7106`].string() // U+7106 <cjk>
	0x8D: [`\u7107`].string() // U+7107 <cjk>
	0x8E: [`\u7108`].string() // U+7108 <cjk>
	0x8F: [`\u710C`].string() // U+710C <cjk>
	0x90: [`\u3DC0`].string() // U+3DC0 <cjk>
	0x91: [`\u712F`].string() // U+712F <cjk>
	0x92: [`\u7131`].string() // U+7131 <cjk>
	0x93: [`\u7150`].string() // U+7150 <cjk>
	0x94: [`\u714A`].string() // U+714A <cjk>
	0x95: [`\u7153`].string() // U+7153 <cjk>
	0x96: [`\u715E`].string() // U+715E <cjk>
	0x97: [`\u3DD4`].string() // U+3DD4 <cjk>
	0x98: [`\u7196`].string() // U+7196 <cjk>
	0x99: [`\u7180`].string() // U+7180 <cjk>
	0x9A: [`\u719B`].string() // U+719B <cjk>
	0x9B: [`\u71A0`].string() // U+71A0 <cjk>
	0x9C: [`\u71A2`].string() // U+71A2 <cjk>
	0x9D: [`\u71AE`].string() // U+71AE <cjk>
	0x9E: [`\u71AF`].string() // U+71AF <cjk>
	0x9F: [`\u71B3`].string() // U+71B3 <cjk>
	0xA0: utf32_to_str(0x243BC) // U+243BC <cjk>
	0xA1: [`\u71CB`].string() // U+71CB <cjk>
	0xA2: [`\u71D3`].string() // U+71D3 <cjk>
	0xA3: [`\u71D9`].string() // U+71D9 <cjk>
	0xA4: [`\u71DC`].string() // U+71DC <cjk>
	0xA5: [`\u7207`].string() // U+7207 <cjk>
	0xA6: [`\u3E05`].string() // U+3E05 <cjk>
	0xA7: [`\uFA49`].string() // U+FA49 CJK COMPATIBILITY IDEOGRAPH-FA49
	0xA8: [`\u722B`].string() // U+722B <cjk>
	0xA9: [`\u7234`].string() // U+7234 <cjk>
	0xAA: [`\u7238`].string() // U+7238 <cjk>
	0xAB: [`\u7239`].string() // U+7239 <cjk>
	0xAC: [`\u4E2C`].string() // U+4E2C <cjk>
	0xAD: [`\u7242`].string() // U+7242 <cjk>
	0xAE: [`\u7253`].string() // U+7253 <cjk>
	0xAF: [`\u7257`].string() // U+7257 <cjk>
	0xB0: [`\u7263`].string() // U+7263 <cjk>
	0xB1: utf32_to_str(0x24629) // U+24629 <cjk>
	0xB2: [`\u726E`].string() // U+726E <cjk>
	0xB3: [`\u726F`].string() // U+726F <cjk>
	0xB4: [`\u7278`].string() // U+7278 <cjk>
	0xB5: [`\u727F`].string() // U+727F <cjk>
	0xB6: [`\u728E`].string() // U+728E <cjk>
	0xB7: utf32_to_str(0x246A5) // U+246A5 <cjk>
	0xB8: [`\u72AD`].string() // U+72AD <cjk>
	0xB9: [`\u72AE`].string() // U+72AE <cjk>
	0xBA: [`\u72B0`].string() // U+72B0 <cjk>
	0xBB: [`\u72B1`].string() // U+72B1 <cjk>
	0xBC: [`\u72C1`].string() // U+72C1 <cjk>
	0xBD: [`\u3E60`].string() // U+3E60 <cjk>
	0xBE: [`\u72CC`].string() // U+72CC <cjk>
	0xBF: [`\u3E66`].string() // U+3E66 <cjk>
	0xC0: [`\u3E68`].string() // U+3E68 <cjk>
	0xC1: [`\u72F3`].string() // U+72F3 <cjk>
	0xC2: [`\u72FA`].string() // U+72FA <cjk>
	0xC3: [`\u7307`].string() // U+7307 <cjk>
	0xC4: [`\u7312`].string() // U+7312 <cjk>
	0xC5: [`\u7318`].string() // U+7318 <cjk>
	0xC6: [`\u7319`].string() // U+7319 <cjk>
	0xC7: [`\u3E83`].string() // U+3E83 <cjk>
	0xC8: [`\u7339`].string() // U+7339 <cjk>
	0xC9: [`\u732C`].string() // U+732C <cjk>
	0xCA: [`\u7331`].string() // U+7331 <cjk>
	0xCB: [`\u7333`].string() // U+7333 <cjk>
	0xCC: [`\u733D`].string() // U+733D <cjk>
	0xCD: [`\u7352`].string() // U+7352 <cjk>
	0xCE: [`\u3E94`].string() // U+3E94 <cjk>
	0xCF: [`\u736B`].string() // U+736B <cjk>
	0xD0: [`\u736C`].string() // U+736C <cjk>
	0xD1: utf32_to_str(0x24896) // U+24896 <cjk>
	0xD2: [`\u736E`].string() // U+736E <cjk>
	0xD3: [`\u736F`].string() // U+736F <cjk>
	0xD4: [`\u7371`].string() // U+7371 <cjk>
	0xD5: [`\u7377`].string() // U+7377 <cjk>
	0xD6: [`\u7381`].string() // U+7381 <cjk>
	0xD7: [`\u7385`].string() // U+7385 <cjk>
	0xD8: [`\u738A`].string() // U+738A <cjk>
	0xD9: [`\u7394`].string() // U+7394 <cjk>
	0xDA: [`\u7398`].string() // U+7398 <cjk>
	0xDB: [`\u739C`].string() // U+739C <cjk>
	0xDC: [`\u739E`].string() // U+739E <cjk>
	0xDD: [`\u73A5`].string() // U+73A5 <cjk>
	0xDE: [`\u73A8`].string() // U+73A8 <cjk>
	0xDF: [`\u73B5`].string() // U+73B5 <cjk>
	0xE0: [`\u73B7`].string() // U+73B7 <cjk>
	0xE1: [`\u73B9`].string() // U+73B9 <cjk>
	0xE2: [`\u73BC`].string() // U+73BC <cjk>
	0xE3: [`\u73BF`].string() // U+73BF <cjk>
	0xE4: [`\u73C5`].string() // U+73C5 <cjk>
	0xE5: [`\u73CB`].string() // U+73CB <cjk>
	0xE6: [`\u73E1`].string() // U+73E1 <cjk>
	0xE7: [`\u73E7`].string() // U+73E7 <cjk>
	0xE8: [`\u73F9`].string() // U+73F9 <cjk>
	0xE9: [`\u7413`].string() // U+7413 <cjk>
	0xEA: [`\u73FA`].string() // U+73FA <cjk>
	0xEB: [`\u7401`].string() // U+7401 <cjk>
	0xEC: [`\u7424`].string() // U+7424 <cjk>
	0xED: [`\u7431`].string() // U+7431 <cjk>
	0xEE: [`\u7439`].string() // U+7439 <cjk>
	0xEF: [`\u7453`].string() // U+7453 <cjk>
	0xF0: [`\u7440`].string() // U+7440 <cjk>
	0xF1: [`\u7443`].string() // U+7443 <cjk>
	0xF2: [`\u744D`].string() // U+744D <cjk>
	0xF3: [`\u7452`].string() // U+7452 <cjk>
	0xF4: [`\u745D`].string() // U+745D <cjk>
	0xF5: [`\u7471`].string() // U+7471 <cjk>
	0xF6: [`\u7481`].string() // U+7481 <cjk>
	0xF7: [`\u7485`].string() // U+7485 <cjk>
	0xF8: [`\u7488`].string() // U+7488 <cjk>
	0xF9: utf32_to_str(0x24A4D) // U+24A4D <cjk>
	0xFA: [`\u7492`].string() // U+7492 <cjk>
	0xFB: [`\u7497`].string() // U+7497 <cjk>
	0xFC: [`\u7499`].string() // U+7499 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x9d = {
	0x40: [`\u621E`].string() // U+621E <cjk>
	0x41: [`\u6221`].string() // U+6221 <cjk>
	0x42: [`\u622A`].string() // U+622A <cjk>
	0x43: [`\u622E`].string() // U+622E <cjk>
	0x44: [`\u6230`].string() // U+6230 <cjk>
	0x45: [`\u6232`].string() // U+6232 <cjk>
	0x46: [`\u6233`].string() // U+6233 <cjk>
	0x47: [`\u6241`].string() // U+6241 <cjk>
	0x48: [`\u624E`].string() // U+624E <cjk>
	0x49: [`\u625E`].string() // U+625E <cjk>
	0x4A: [`\u6263`].string() // U+6263 <cjk>
	0x4B: [`\u625B`].string() // U+625B <cjk>
	0x4C: [`\u6260`].string() // U+6260 <cjk>
	0x4D: [`\u6268`].string() // U+6268 <cjk>
	0x4E: [`\u627C`].string() // U+627C <cjk>
	0x4F: [`\u6282`].string() // U+6282 <cjk>
	0x50: [`\u6289`].string() // U+6289 <cjk>
	0x51: [`\u627E`].string() // U+627E <cjk>
	0x52: [`\u6292`].string() // U+6292 <cjk>
	0x53: [`\u6293`].string() // U+6293 <cjk>
	0x54: [`\u6296`].string() // U+6296 <cjk>
	0x55: [`\u62D4`].string() // U+62D4 <cjk>
	0x56: [`\u6283`].string() // U+6283 <cjk>
	0x57: [`\u6294`].string() // U+6294 <cjk>
	0x58: [`\u62D7`].string() // U+62D7 <cjk>
	0x59: [`\u62D1`].string() // U+62D1 <cjk>
	0x5A: [`\u62BB`].string() // U+62BB <cjk>
	0x5B: [`\u62CF`].string() // U+62CF <cjk>
	0x5C: [`\u62FF`].string() // U+62FF <cjk>
	0x5D: [`\u62C6`].string() // U+62C6 <cjk>
	0x5E: [`\u64D4`].string() // U+64D4 <cjk>
	0x5F: [`\u62C8`].string() // U+62C8 <cjk>
	0x60: [`\u62DC`].string() // U+62DC <cjk>
	0x61: [`\u62CC`].string() // U+62CC <cjk>
	0x62: [`\u62CA`].string() // U+62CA <cjk>
	0x63: [`\u62C2`].string() // U+62C2 <cjk>
	0x64: [`\u62C7`].string() // U+62C7 <cjk>
	0x65: [`\u629B`].string() // U+629B <cjk>
	0x66: [`\u62C9`].string() // U+62C9 <cjk>
	0x67: [`\u630C`].string() // U+630C <cjk>
	0x68: [`\u62EE`].string() // U+62EE <cjk>
	0x69: [`\u62F1`].string() // U+62F1 <cjk>
	0x6A: [`\u6327`].string() // U+6327 <cjk>
	0x6B: [`\u6302`].string() // U+6302 <cjk>
	0x6C: [`\u6308`].string() // U+6308 <cjk>
	0x6D: [`\u62EF`].string() // U+62EF <cjk>
	0x6E: [`\u62F5`].string() // U+62F5 <cjk>
	0x6F: [`\u6350`].string() // U+6350 <cjk>
	0x70: [`\u633E`].string() // U+633E <cjk>
	0x71: [`\u634D`].string() // U+634D <cjk>
	0x72: [`\u641C`].string() // U+641C <cjk>
	0x73: [`\u634F`].string() // U+634F <cjk>
	0x74: [`\u6396`].string() // U+6396 <cjk>
	0x75: [`\u638E`].string() // U+638E <cjk>
	0x76: [`\u6380`].string() // U+6380 <cjk>
	0x77: [`\u63AB`].string() // U+63AB <cjk>
	0x78: [`\u6376`].string() // U+6376 <cjk>
	0x79: [`\u63A3`].string() // U+63A3 <cjk>
	0x7A: [`\u638F`].string() // U+638F <cjk>
	0x7B: [`\u6389`].string() // U+6389 <cjk>
	0x7C: [`\u639F`].string() // U+639F <cjk>
	0x7D: [`\u63B5`].string() // U+63B5 <cjk>
	0x7E: [`\u636B`].string() // U+636B <cjk>
	0x80: [`\u6369`].string() // U+6369 <cjk>
	0x81: [`\u63BE`].string() // U+63BE <cjk>
	0x82: [`\u63E9`].string() // U+63E9 <cjk>
	0x83: [`\u63C0`].string() // U+63C0 <cjk>
	0x84: [`\u63C6`].string() // U+63C6 <cjk>
	0x85: [`\u63E3`].string() // U+63E3 <cjk>
	0x86: [`\u63C9`].string() // U+63C9 <cjk>
	0x87: [`\u63D2`].string() // U+63D2 <cjk>
	0x88: [`\u63F6`].string() // U+63F6 <cjk>
	0x89: [`\u63C4`].string() // U+63C4 <cjk>
	0x8A: [`\u6416`].string() // U+6416 <cjk>
	0x8B: [`\u6434`].string() // U+6434 <cjk>
	0x8C: [`\u6406`].string() // U+6406 <cjk>
	0x8D: [`\u6413`].string() // U+6413 <cjk>
	0x8E: [`\u6426`].string() // U+6426 <cjk>
	0x8F: [`\u6436`].string() // U+6436 <cjk>
	0x90: [`\u651D`].string() // U+651D <cjk>
	0x91: [`\u6417`].string() // U+6417 <cjk>
	0x92: [`\u6428`].string() // U+6428 <cjk>
	0x93: [`\u640F`].string() // U+640F <cjk>
	0x94: [`\u6467`].string() // U+6467 <cjk>
	0x95: [`\u646F`].string() // U+646F <cjk>
	0x96: [`\u6476`].string() // U+6476 <cjk>
	0x97: [`\u644E`].string() // U+644E <cjk>
	0x98: [`\u652A`].string() // U+652A <cjk>
	0x99: [`\u6495`].string() // U+6495 <cjk>
	0x9A: [`\u6493`].string() // U+6493 <cjk>
	0x9B: [`\u64A5`].string() // U+64A5 <cjk>
	0x9C: [`\u64A9`].string() // U+64A9 <cjk>
	0x9D: [`\u6488`].string() // U+6488 <cjk>
	0x9E: [`\u64BC`].string() // U+64BC <cjk>
	0x9F: [`\u64DA`].string() // U+64DA <cjk>
	0xA0: [`\u64D2`].string() // U+64D2 <cjk>
	0xA1: [`\u64C5`].string() // U+64C5 <cjk>
	0xA2: [`\u64C7`].string() // U+64C7 <cjk>
	0xA3: [`\u64BB`].string() // U+64BB <cjk>
	0xA4: [`\u64D8`].string() // U+64D8 <cjk>
	0xA5: [`\u64C2`].string() // U+64C2 <cjk>
	0xA6: [`\u64F1`].string() // U+64F1 <cjk>
	0xA7: [`\u64E7`].string() // U+64E7 <cjk>
	0xA8: [`\u8209`].string() // U+8209 <cjk>
	0xA9: [`\u64E0`].string() // U+64E0 <cjk>
	0xAA: [`\u64E1`].string() // U+64E1 <cjk>
	0xAB: [`\u62AC`].string() // U+62AC <cjk>
	0xAC: [`\u64E3`].string() // U+64E3 <cjk>
	0xAD: [`\u64EF`].string() // U+64EF <cjk>
	0xAE: [`\u652C`].string() // U+652C <cjk>
	0xAF: [`\u64F6`].string() // U+64F6 <cjk>
	0xB0: [`\u64F4`].string() // U+64F4 <cjk>
	0xB1: [`\u64F2`].string() // U+64F2 <cjk>
	0xB2: [`\u64FA`].string() // U+64FA <cjk>
	0xB3: [`\u6500`].string() // U+6500 <cjk>
	0xB4: [`\u64FD`].string() // U+64FD <cjk>
	0xB5: [`\u6518`].string() // U+6518 <cjk>
	0xB6: [`\u651C`].string() // U+651C <cjk>
	0xB7: [`\u6505`].string() // U+6505 <cjk>
	0xB8: [`\u6524`].string() // U+6524 <cjk>
	0xB9: [`\u6523`].string() // U+6523 <cjk>
	0xBA: [`\u652B`].string() // U+652B <cjk>
	0xBB: [`\u6534`].string() // U+6534 <cjk>
	0xBC: [`\u6535`].string() // U+6535 <cjk>
	0xBD: [`\u6537`].string() // U+6537 <cjk>
	0xBE: [`\u6536`].string() // U+6536 <cjk>
	0xBF: [`\u6538`].string() // U+6538 <cjk>
	0xC0: [`\u754B`].string() // U+754B <cjk>
	0xC1: [`\u6548`].string() // U+6548 <cjk>
	0xC2: [`\u6556`].string() // U+6556 <cjk>
	0xC3: [`\u6555`].string() // U+6555 <cjk>
	0xC4: [`\u654D`].string() // U+654D <cjk>
	0xC5: [`\u6558`].string() // U+6558 <cjk>
	0xC6: [`\u655E`].string() // U+655E <cjk>
	0xC7: [`\u655D`].string() // U+655D <cjk>
	0xC8: [`\u6572`].string() // U+6572 <cjk>
	0xC9: [`\u6578`].string() // U+6578 <cjk>
	0xCA: [`\u6582`].string() // U+6582 <cjk>
	0xCB: [`\u6583`].string() // U+6583 <cjk>
	0xCC: [`\u8B8A`].string() // U+8B8A <cjk>
	0xCD: [`\u659B`].string() // U+659B <cjk>
	0xCE: [`\u659F`].string() // U+659F <cjk>
	0xCF: [`\u65AB`].string() // U+65AB <cjk>
	0xD0: [`\u65B7`].string() // U+65B7 <cjk>
	0xD1: [`\u65C3`].string() // U+65C3 <cjk>
	0xD2: [`\u65C6`].string() // U+65C6 <cjk>
	0xD3: [`\u65C1`].string() // U+65C1 <cjk>
	0xD4: [`\u65C4`].string() // U+65C4 <cjk>
	0xD5: [`\u65CC`].string() // U+65CC <cjk>
	0xD6: [`\u65D2`].string() // U+65D2 <cjk>
	0xD7: [`\u65DB`].string() // U+65DB <cjk>
	0xD8: [`\u65D9`].string() // U+65D9 <cjk>
	0xD9: [`\u65E0`].string() // U+65E0 <cjk>
	0xDA: [`\u65E1`].string() // U+65E1 <cjk>
	0xDB: [`\u65F1`].string() // U+65F1 <cjk>
	0xDC: [`\u6772`].string() // U+6772 <cjk>
	0xDD: [`\u660A`].string() // U+660A <cjk>
	0xDE: [`\u6603`].string() // U+6603 <cjk>
	0xDF: [`\u65FB`].string() // U+65FB <cjk>
	0xE0: [`\u6773`].string() // U+6773 <cjk>
	0xE1: [`\u6635`].string() // U+6635 <cjk>
	0xE2: [`\u6636`].string() // U+6636 <cjk>
	0xE3: [`\u6634`].string() // U+6634 <cjk>
	0xE4: [`\u661C`].string() // U+661C <cjk>
	0xE5: [`\u664F`].string() // U+664F <cjk>
	0xE6: [`\u6644`].string() // U+6644 <cjk>
	0xE7: [`\u6649`].string() // U+6649 <cjk>
	0xE8: [`\u6641`].string() // U+6641 <cjk>
	0xE9: [`\u665E`].string() // U+665E <cjk>
	0xEA: [`\u665D`].string() // U+665D <cjk>
	0xEB: [`\u6664`].string() // U+6664 <cjk>
	0xEC: [`\u6667`].string() // U+6667 <cjk>
	0xED: [`\u6668`].string() // U+6668 <cjk>
	0xEE: [`\u665F`].string() // U+665F <cjk>
	0xEF: [`\u6662`].string() // U+6662 <cjk>
	0xF0: [`\u6670`].string() // U+6670 <cjk>
	0xF1: [`\u6683`].string() // U+6683 <cjk>
	0xF2: [`\u6688`].string() // U+6688 <cjk>
	0xF3: [`\u668E`].string() // U+668E <cjk>
	0xF4: [`\u6689`].string() // U+6689 <cjk>
	0xF5: [`\u6684`].string() // U+6684 <cjk>
	0xF6: [`\u6698`].string() // U+6698 <cjk>
	0xF7: [`\u669D`].string() // U+669D <cjk>
	0xF8: [`\u66C1`].string() // U+66C1 <cjk>
	0xF9: [`\u66B9`].string() // U+66B9 <cjk>
	0xFA: [`\u66C9`].string() // U+66C9 <cjk>
	0xFB: [`\u66BE`].string() // U+66BE <cjk>
	0xFC: [`\u66BC`].string() // U+66BC <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xfa = {
	0x40: [`\u8C57`].string() // U+8C57 <cjk>
	0x41: [`\u8C69`].string() // U+8C69 <cjk>
	0x42: [`\u8C6D`].string() // U+8C6D <cjk>
	0x43: [`\u8C73`].string() // U+8C73 <cjk>
	0x44: utf32_to_str(0x27CB8) // U+27CB8 <cjk>
	0x45: [`\u8C93`].string() // U+8C93 <cjk>
	0x46: [`\u8C92`].string() // U+8C92 <cjk>
	0x47: [`\u8C99`].string() // U+8C99 <cjk>
	0x48: [`\u4764`].string() // U+4764 <cjk>
	0x49: [`\u8C9B`].string() // U+8C9B <cjk>
	0x4A: [`\u8CA4`].string() // U+8CA4 <cjk>
	0x4B: [`\u8CD6`].string() // U+8CD6 <cjk>
	0x4C: [`\u8CD5`].string() // U+8CD5 <cjk>
	0x4D: [`\u8CD9`].string() // U+8CD9 <cjk>
	0x4E: utf32_to_str(0x27DA0) // U+27DA0 <cjk>
	0x4F: [`\u8CF0`].string() // U+8CF0 <cjk>
	0x50: [`\u8CF1`].string() // U+8CF1 <cjk>
	0x51: utf32_to_str(0x27E10) // U+27E10 <cjk>
	0x52: [`\u8D09`].string() // U+8D09 <cjk>
	0x53: [`\u8D0E`].string() // U+8D0E <cjk>
	0x54: [`\u8D6C`].string() // U+8D6C <cjk>
	0x55: [`\u8D84`].string() // U+8D84 <cjk>
	0x56: [`\u8D95`].string() // U+8D95 <cjk>
	0x57: [`\u8DA6`].string() // U+8DA6 <cjk>
	0x58: utf32_to_str(0x27FB7) // U+27FB7 <cjk>
	0x59: [`\u8DC6`].string() // U+8DC6 <cjk>
	0x5A: [`\u8DC8`].string() // U+8DC8 <cjk>
	0x5B: [`\u8DD9`].string() // U+8DD9 <cjk>
	0x5C: [`\u8DEC`].string() // U+8DEC <cjk>
	0x5D: [`\u8E0C`].string() // U+8E0C <cjk>
	0x5E: [`\u47FD`].string() // U+47FD <cjk>
	0x5F: [`\u8DFD`].string() // U+8DFD <cjk>
	0x60: [`\u8E06`].string() // U+8E06 <cjk>
	0x61: utf32_to_str(0x2808A) // U+2808A <cjk>
	0x62: [`\u8E14`].string() // U+8E14 <cjk>
	0x63: [`\u8E16`].string() // U+8E16 <cjk>
	0x64: [`\u8E21`].string() // U+8E21 <cjk>
	0x65: [`\u8E22`].string() // U+8E22 <cjk>
	0x66: [`\u8E27`].string() // U+8E27 <cjk>
	0x67: utf32_to_str(0x280BB) // U+280BB <cjk>
	0x68: [`\u4816`].string() // U+4816 <cjk>
	0x69: [`\u8E36`].string() // U+8E36 <cjk>
	0x6A: [`\u8E39`].string() // U+8E39 <cjk>
	0x6B: [`\u8E4B`].string() // U+8E4B <cjk>
	0x6C: [`\u8E54`].string() // U+8E54 <cjk>
	0x6D: [`\u8E62`].string() // U+8E62 <cjk>
	0x6E: [`\u8E6C`].string() // U+8E6C <cjk>
	0x6F: [`\u8E6D`].string() // U+8E6D <cjk>
	0x70: [`\u8E6F`].string() // U+8E6F <cjk>
	0x71: [`\u8E98`].string() // U+8E98 <cjk>
	0x72: [`\u8E9E`].string() // U+8E9E <cjk>
	0x73: [`\u8EAE`].string() // U+8EAE <cjk>
	0x74: [`\u8EB3`].string() // U+8EB3 <cjk>
	0x75: [`\u8EB5`].string() // U+8EB5 <cjk>
	0x76: [`\u8EB6`].string() // U+8EB6 <cjk>
	0x77: [`\u8EBB`].string() // U+8EBB <cjk>
	0x78: utf32_to_str(0x28282) // U+28282 <cjk>
	0x79: [`\u8ED1`].string() // U+8ED1 <cjk>
	0x7A: [`\u8ED4`].string() // U+8ED4 <cjk>
	0x7B: [`\u484E`].string() // U+484E <cjk>
	0x7C: [`\u8EF9`].string() // U+8EF9 <cjk>
	0x7D: utf32_to_str(0x282F3) // U+282F3 <cjk>
	0x7E: [`\u8F00`].string() // U+8F00 <cjk>
	0x80: [`\u8F08`].string() // U+8F08 <cjk>
	0x81: [`\u8F17`].string() // U+8F17 <cjk>
	0x82: [`\u8F2B`].string() // U+8F2B <cjk>
	0x83: [`\u8F40`].string() // U+8F40 <cjk>
	0x84: [`\u8F4A`].string() // U+8F4A <cjk>
	0x85: [`\u8F58`].string() // U+8F58 <cjk>
	0x86: utf32_to_str(0x2840C) // U+2840C <cjk>
	0x87: [`\u8FA4`].string() // U+8FA4 <cjk>
	0x88: [`\u8FB4`].string() // U+8FB4 <cjk>
	0x89: [`\uFA66`].string() // U+FA66 CJK COMPATIBILITY IDEOGRAPH-FA66
	0x8A: [`\u8FB6`].string() // U+8FB6 <cjk>
	0x8B: utf32_to_str(0x28455) // U+28455 <cjk>
	0x8C: [`\u8FC1`].string() // U+8FC1 <cjk>
	0x8D: [`\u8FC6`].string() // U+8FC6 <cjk>
	0x8E: [`\uFA24`].string() // U+FA24 CJK COMPATIBILITY IDEOGRAPH-FA24
	0x8F: [`\u8FCA`].string() // U+8FCA <cjk>
	0x90: [`\u8FCD`].string() // U+8FCD <cjk>
	0x91: [`\u8FD3`].string() // U+8FD3 <cjk>
	0x92: [`\u8FD5`].string() // U+8FD5 <cjk>
	0x93: [`\u8FE0`].string() // U+8FE0 <cjk>
	0x94: [`\u8FF1`].string() // U+8FF1 <cjk>
	0x95: [`\u8FF5`].string() // U+8FF5 <cjk>
	0x96: [`\u8FFB`].string() // U+8FFB <cjk>
	0x97: [`\u9002`].string() // U+9002 <cjk>
	0x98: [`\u900C`].string() // U+900C <cjk>
	0x99: [`\u9037`].string() // U+9037 <cjk>
	0x9A: utf32_to_str(0x2856B) // U+2856B <cjk>
	0x9B: [`\u9043`].string() // U+9043 <cjk>
	0x9C: [`\u9044`].string() // U+9044 <cjk>
	0x9D: [`\u905D`].string() // U+905D <cjk>
	0x9E: utf32_to_str(0x285C8) // U+285C8 <cjk>
	0x9F: utf32_to_str(0x285C9) // U+285C9 <cjk>
	0xA0: [`\u9085`].string() // U+9085 <cjk>
	0xA1: [`\u908C`].string() // U+908C <cjk>
	0xA2: [`\u9090`].string() // U+9090 <cjk>
	0xA3: [`\u961D`].string() // U+961D <cjk>
	0xA4: [`\u90A1`].string() // U+90A1 <cjk>
	0xA5: [`\u48B5`].string() // U+48B5 <cjk>
	0xA6: [`\u90B0`].string() // U+90B0 <cjk>
	0xA7: [`\u90B6`].string() // U+90B6 <cjk>
	0xA8: [`\u90C3`].string() // U+90C3 <cjk>
	0xA9: [`\u90C8`].string() // U+90C8 <cjk>
	0xAA: utf32_to_str(0x286D7) // U+286D7 <cjk>
	0xAB: [`\u90DC`].string() // U+90DC <cjk>
	0xAC: [`\u90DF`].string() // U+90DF <cjk>
	0xAD: utf32_to_str(0x286FA) // U+286FA <cjk>
	0xAE: [`\u90F6`].string() // U+90F6 <cjk>
	0xAF: [`\u90F2`].string() // U+90F2 <cjk>
	0xB0: [`\u9100`].string() // U+9100 <cjk>
	0xB1: [`\u90EB`].string() // U+90EB <cjk>
	0xB2: [`\u90FE`].string() // U+90FE <cjk>
	0xB3: [`\u90FF`].string() // U+90FF <cjk>
	0xB4: [`\u9104`].string() // U+9104 <cjk>
	0xB5: [`\u9106`].string() // U+9106 <cjk>
	0xB6: [`\u9118`].string() // U+9118 <cjk>
	0xB7: [`\u911C`].string() // U+911C <cjk>
	0xB8: [`\u911E`].string() // U+911E <cjk>
	0xB9: [`\u9137`].string() // U+9137 <cjk>
	0xBA: [`\u9139`].string() // U+9139 <cjk>
	0xBB: [`\u913A`].string() // U+913A <cjk>
	0xBC: [`\u9146`].string() // U+9146 <cjk>
	0xBD: [`\u9147`].string() // U+9147 <cjk>
	0xBE: [`\u9157`].string() // U+9157 <cjk>
	0xBF: [`\u9159`].string() // U+9159 <cjk>
	0xC0: [`\u9161`].string() // U+9161 <cjk>
	0xC1: [`\u9164`].string() // U+9164 <cjk>
	0xC2: [`\u9174`].string() // U+9174 <cjk>
	0xC3: [`\u9179`].string() // U+9179 <cjk>
	0xC4: [`\u9185`].string() // U+9185 <cjk>
	0xC5: [`\u918E`].string() // U+918E <cjk>
	0xC6: [`\u91A8`].string() // U+91A8 <cjk>
	0xC7: [`\u91AE`].string() // U+91AE <cjk>
	0xC8: [`\u91B3`].string() // U+91B3 <cjk>
	0xC9: [`\u91B6`].string() // U+91B6 <cjk>
	0xCA: [`\u91C3`].string() // U+91C3 <cjk>
	0xCB: [`\u91C4`].string() // U+91C4 <cjk>
	0xCC: [`\u91DA`].string() // U+91DA <cjk>
	0xCD: utf32_to_str(0x28949) // U+28949 <cjk>
	0xCE: utf32_to_str(0x28946) // U+28946 <cjk>
	0xCF: [`\u91EC`].string() // U+91EC <cjk>
	0xD0: [`\u91EE`].string() // U+91EE <cjk>
	0xD1: [`\u9201`].string() // U+9201 <cjk>
	0xD2: [`\u920A`].string() // U+920A <cjk>
	0xD3: [`\u9216`].string() // U+9216 <cjk>
	0xD4: [`\u9217`].string() // U+9217 <cjk>
	0xD5: utf32_to_str(0x2896B) // U+2896B <cjk>
	0xD6: [`\u9233`].string() // U+9233 <cjk>
	0xD7: [`\u9242`].string() // U+9242 <cjk>
	0xD8: [`\u9247`].string() // U+9247 <cjk>
	0xD9: [`\u924A`].string() // U+924A <cjk>
	0xDA: [`\u924E`].string() // U+924E <cjk>
	0xDB: [`\u9251`].string() // U+9251 <cjk>
	0xDC: [`\u9256`].string() // U+9256 <cjk>
	0xDD: [`\u9259`].string() // U+9259 <cjk>
	0xDE: [`\u9260`].string() // U+9260 <cjk>
	0xDF: [`\u9261`].string() // U+9261 <cjk>
	0xE0: [`\u9265`].string() // U+9265 <cjk>
	0xE1: [`\u9267`].string() // U+9267 <cjk>
	0xE2: [`\u9268`].string() // U+9268 <cjk>
	0xE3: utf32_to_str(0x28987) // U+28987 <cjk>
	0xE4: utf32_to_str(0x28988) // U+28988 <cjk>
	0xE5: [`\u927C`].string() // U+927C <cjk>
	0xE6: [`\u927D`].string() // U+927D <cjk>
	0xE7: [`\u927F`].string() // U+927F <cjk>
	0xE8: [`\u9289`].string() // U+9289 <cjk>
	0xE9: [`\u928D`].string() // U+928D <cjk>
	0xEA: [`\u9297`].string() // U+9297 <cjk>
	0xEB: [`\u9299`].string() // U+9299 <cjk>
	0xEC: [`\u929F`].string() // U+929F <cjk>
	0xED: [`\u92A7`].string() // U+92A7 <cjk>
	0xEE: [`\u92AB`].string() // U+92AB <cjk>
	0xEF: utf32_to_str(0x289BA) // U+289BA <cjk>
	0xF0: utf32_to_str(0x289BB) // U+289BB <cjk>
	0xF1: [`\u92B2`].string() // U+92B2 <cjk>
	0xF2: [`\u92BF`].string() // U+92BF <cjk>
	0xF3: [`\u92C0`].string() // U+92C0 <cjk>
	0xF4: [`\u92C6`].string() // U+92C6 <cjk>
	0xF5: [`\u92CE`].string() // U+92CE <cjk>
	0xF6: [`\u92D0`].string() // U+92D0 <cjk>
	0xF7: [`\u92D7`].string() // U+92D7 <cjk>
	0xF8: [`\u92D9`].string() // U+92D9 <cjk>
	0xF9: [`\u92E5`].string() // U+92E5 <cjk>
	0xFA: [`\u92E7`].string() // U+92E7 <cjk>
	0xFB: [`\u9311`].string() // U+9311 <cjk>
	0xFC: utf32_to_str(0x28A1E) // U+28A1E <cjk>
}

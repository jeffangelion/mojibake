module mojibake

const jis_x_0213_doublebyte_0xec = {
	0x40: [`\u6EC7`].string() // U+6EC7 <cjk>
	0x41: [`\u6ECE`].string() // U+6ECE <cjk>
	0x42: [`\u6F10`].string() // U+6F10 <cjk>
	0x43: [`\u6F1A`].string() // U+6F1A <cjk>
	0x44: [`\uFA47`].string() // U+FA47 CJK COMPATIBILITY IDEOGRAPH-FA47
	0x45: [`\u6F2A`].string() // U+6F2A <cjk>
	0x46: [`\u6F2F`].string() // U+6F2F <cjk>
	0x47: [`\u6F33`].string() // U+6F33 <cjk>
	0x48: [`\u6F51`].string() // U+6F51 <cjk>
	0x49: [`\u6F59`].string() // U+6F59 <cjk>
	0x4A: [`\u6F5E`].string() // U+6F5E <cjk>
	0x4B: [`\u6F61`].string() // U+6F61 <cjk>
	0x4C: [`\u6F62`].string() // U+6F62 <cjk>
	0x4D: [`\u6F7E`].string() // U+6F7E <cjk>
	0x4E: [`\u6F88`].string() // U+6F88 <cjk>
	0x4F: [`\u6F8C`].string() // U+6F8C <cjk>
	0x50: [`\u6F8D`].string() // U+6F8D <cjk>
	0x51: [`\u6F94`].string() // U+6F94 <cjk>
	0x52: [`\u6FA0`].string() // U+6FA0 <cjk>
	0x53: [`\u6FA7`].string() // U+6FA7 <cjk>
	0x54: [`\u6FB6`].string() // U+6FB6 <cjk>
	0x55: [`\u6FBC`].string() // U+6FBC <cjk>
	0x56: [`\u6FC7`].string() // U+6FC7 <cjk>
	0x57: [`\u6FCA`].string() // U+6FCA <cjk>
	0x58: [`\u6FF9`].string() // U+6FF9 <cjk>
	0x59: [`\u6FF0`].string() // U+6FF0 <cjk>
	0x5A: [`\u6FF5`].string() // U+6FF5 <cjk>
	0x5B: [`\u7005`].string() // U+7005 <cjk>
	0x5C: [`\u7006`].string() // U+7006 <cjk>
	0x5D: [`\u7028`].string() // U+7028 <cjk>
	0x5E: [`\u704A`].string() // U+704A <cjk>
	0x5F: [`\u705D`].string() // U+705D <cjk>
	0x60: [`\u705E`].string() // U+705E <cjk>
	0x61: [`\u704E`].string() // U+704E <cjk>
	0x62: [`\u7064`].string() // U+7064 <cjk>
	0x63: [`\u7075`].string() // U+7075 <cjk>
	0x64: [`\u7085`].string() // U+7085 <cjk>
	0x65: [`\u70A4`].string() // U+70A4 <cjk>
	0x66: [`\u70AB`].string() // U+70AB <cjk>
	0x67: [`\u70B7`].string() // U+70B7 <cjk>
	0x68: [`\u70D4`].string() // U+70D4 <cjk>
	0x69: [`\u70D8`].string() // U+70D8 <cjk>
	0x6A: [`\u70E4`].string() // U+70E4 <cjk>
	0x6B: [`\u710F`].string() // U+710F <cjk>
	0x6C: [`\u712B`].string() // U+712B <cjk>
	0x6D: [`\u711E`].string() // U+711E <cjk>
	0x6E: [`\u7120`].string() // U+7120 <cjk>
	0x6F: [`\u712E`].string() // U+712E <cjk>
	0x70: [`\u7130`].string() // U+7130 <cjk>
	0x71: [`\u7146`].string() // U+7146 <cjk>
	0x72: [`\u7147`].string() // U+7147 <cjk>
	0x73: [`\u7151`].string() // U+7151 <cjk>
	0x74: [`\uFA48`].string() // U+FA48 CJK COMPATIBILITY IDEOGRAPH-FA48
	0x75: [`\u7152`].string() // U+7152 <cjk>
	0x76: [`\u715C`].string() // U+715C <cjk>
	0x77: [`\u7160`].string() // U+7160 <cjk>
	0x78: [`\u7168`].string() // U+7168 <cjk>
	0x79: [`\uFA15`].string() // U+FA15 CJK COMPATIBILITY IDEOGRAPH-FA15
	0x7A: [`\u7185`].string() // U+7185 <cjk>
	0x7B: [`\u7187`].string() // U+7187 <cjk>
	0x7C: [`\u7192`].string() // U+7192 <cjk>
	0x7D: [`\u71C1`].string() // U+71C1 <cjk>
	0x7E: [`\u71BA`].string() // U+71BA <cjk>
	0x80: [`\u71C4`].string() // U+71C4 <cjk>
	0x81: [`\u71FE`].string() // U+71FE <cjk>
	0x82: [`\u7200`].string() // U+7200 <cjk>
	0x83: [`\u7215`].string() // U+7215 <cjk>
	0x84: [`\u7255`].string() // U+7255 <cjk>
	0x85: [`\u7256`].string() // U+7256 <cjk>
	0x86: [`\u3E3F`].string() // U+3E3F <cjk>
	0x87: [`\u728D`].string() // U+728D <cjk>
	0x88: [`\u729B`].string() // U+729B <cjk>
	0x89: [`\u72BE`].string() // U+72BE <cjk>
	0x8A: [`\u72C0`].string() // U+72C0 <cjk>
	0x8B: [`\u72FB`].string() // U+72FB <cjk>
	0x8C: utf32_to_str(0x247F1) // U+247F1 <cjk>
	0x8D: [`\u7327`].string() // U+7327 <cjk>
	0x8E: [`\u7328`].string() // U+7328 <cjk>
	0x8F: [`\uFA16`].string() // U+FA16 CJK COMPATIBILITY IDEOGRAPH-FA16
	0x90: [`\u7350`].string() // U+7350 <cjk>
	0x91: [`\u7366`].string() // U+7366 <cjk>
	0x92: [`\u737C`].string() // U+737C <cjk>
	0x93: [`\u7395`].string() // U+7395 <cjk>
	0x94: [`\u739F`].string() // U+739F <cjk>
	0x95: [`\u73A0`].string() // U+73A0 <cjk>
	0x96: [`\u73A2`].string() // U+73A2 <cjk>
	0x97: [`\u73A6`].string() // U+73A6 <cjk>
	0x98: [`\u73AB`].string() // U+73AB <cjk>
	0x99: [`\u73C9`].string() // U+73C9 <cjk>
	0x9A: [`\u73CF`].string() // U+73CF <cjk>
	0x9B: [`\u73D6`].string() // U+73D6 <cjk>
	0x9C: [`\u73D9`].string() // U+73D9 <cjk>
	0x9D: [`\u73E3`].string() // U+73E3 <cjk>
	0x9E: [`\u73E9`].string() // U+73E9 <cjk>
	0x9F: [`\u7407`].string() // U+7407 <cjk>
	0xA0: [`\u740A`].string() // U+740A <cjk>
	0xA1: [`\u741A`].string() // U+741A <cjk>
	0xA2: [`\u741B`].string() // U+741B <cjk>
	0xA3: [`\uFA4A`].string() // U+FA4A CJK COMPATIBILITY IDEOGRAPH-FA4A
	0xA4: [`\u7426`].string() // U+7426 <cjk>
	0xA5: [`\u7428`].string() // U+7428 <cjk>
	0xA6: [`\u742A`].string() // U+742A <cjk>
	0xA7: [`\u742B`].string() // U+742B <cjk>
	0xA8: [`\u742C`].string() // U+742C <cjk>
	0xA9: [`\u742E`].string() // U+742E <cjk>
	0xAA: [`\u742F`].string() // U+742F <cjk>
	0xAB: [`\u7430`].string() // U+7430 <cjk>
	0xAC: [`\u7444`].string() // U+7444 <cjk>
	0xAD: [`\u7446`].string() // U+7446 <cjk>
	0xAE: [`\u7447`].string() // U+7447 <cjk>
	0xAF: [`\u744B`].string() // U+744B <cjk>
	0xB0: [`\u7457`].string() // U+7457 <cjk>
	0xB1: [`\u7462`].string() // U+7462 <cjk>
	0xB2: [`\u746B`].string() // U+746B <cjk>
	0xB3: [`\u746D`].string() // U+746D <cjk>
	0xB4: [`\u7486`].string() // U+7486 <cjk>
	0xB5: [`\u7487`].string() // U+7487 <cjk>
	0xB6: [`\u7489`].string() // U+7489 <cjk>
	0xB7: [`\u7498`].string() // U+7498 <cjk>
	0xB8: [`\u749C`].string() // U+749C <cjk>
	0xB9: [`\u749F`].string() // U+749F <cjk>
	0xBA: [`\u74A3`].string() // U+74A3 <cjk>
	0xBB: [`\u7490`].string() // U+7490 <cjk>
	0xBC: [`\u74A6`].string() // U+74A6 <cjk>
	0xBD: [`\u74A8`].string() // U+74A8 <cjk>
	0xBE: [`\u74A9`].string() // U+74A9 <cjk>
	0xBF: [`\u74B5`].string() // U+74B5 <cjk>
	0xC0: [`\u74BF`].string() // U+74BF <cjk>
	0xC1: [`\u74C8`].string() // U+74C8 <cjk>
	0xC2: [`\u74C9`].string() // U+74C9 <cjk>
	0xC3: [`\u74DA`].string() // U+74DA <cjk>
	0xC4: [`\u74FF`].string() // U+74FF <cjk>
	0xC5: [`\u7501`].string() // U+7501 <cjk>
	0xC6: [`\u7517`].string() // U+7517 <cjk>
	0xC7: [`\u752F`].string() // U+752F <cjk>
	0xC8: [`\u756F`].string() // U+756F <cjk>
	0xC9: [`\u7579`].string() // U+7579 <cjk>
	0xCA: [`\u7592`].string() // U+7592 <cjk>
	0xCB: [`\u3F72`].string() // U+3F72 <cjk>
	0xCC: [`\u75CE`].string() // U+75CE <cjk>
	0xCD: [`\u75E4`].string() // U+75E4 <cjk>
	0xCE: [`\u7600`].string() // U+7600 <cjk>
	0xCF: [`\u7602`].string() // U+7602 <cjk>
	0xD0: [`\u7608`].string() // U+7608 <cjk>
	0xD1: [`\u7615`].string() // U+7615 <cjk>
	0xD2: [`\u7616`].string() // U+7616 <cjk>
	0xD3: [`\u7619`].string() // U+7619 <cjk>
	0xD4: [`\u761E`].string() // U+761E <cjk>
	0xD5: [`\u762D`].string() // U+762D <cjk>
	0xD6: [`\u7635`].string() // U+7635 <cjk>
	0xD7: [`\u7643`].string() // U+7643 <cjk>
	0xD8: [`\u764B`].string() // U+764B <cjk>
	0xD9: [`\u7664`].string() // U+7664 <cjk>
	0xDA: [`\u7665`].string() // U+7665 <cjk>
	0xDB: [`\u766D`].string() // U+766D <cjk>
	0xDC: [`\u766F`].string() // U+766F <cjk>
	0xDD: [`\u7671`].string() // U+7671 <cjk>
	0xDE: [`\u7681`].string() // U+7681 <cjk>
	0xDF: [`\u769B`].string() // U+769B <cjk>
	0xE0: [`\u769D`].string() // U+769D <cjk>
	0xE1: [`\u769E`].string() // U+769E <cjk>
	0xE2: [`\u76A6`].string() // U+76A6 <cjk>
	0xE3: [`\u76AA`].string() // U+76AA <cjk>
	0xE4: [`\u76B6`].string() // U+76B6 <cjk>
	0xE5: [`\u76C5`].string() // U+76C5 <cjk>
	0xE6: [`\u76CC`].string() // U+76CC <cjk>
	0xE7: [`\u76CE`].string() // U+76CE <cjk>
	0xE8: [`\u76D4`].string() // U+76D4 <cjk>
	0xE9: [`\u76E6`].string() // U+76E6 <cjk>
	0xEA: [`\u76F1`].string() // U+76F1 <cjk>
	0xEB: [`\u76FC`].string() // U+76FC <cjk>
	0xEC: [`\u770A`].string() // U+770A <cjk>
	0xED: [`\u7719`].string() // U+7719 <cjk>
	0xEE: [`\u7734`].string() // U+7734 <cjk>
	0xEF: [`\u7736`].string() // U+7736 <cjk>
	0xF0: [`\u7746`].string() // U+7746 <cjk>
	0xF1: [`\u774D`].string() // U+774D <cjk>
	0xF2: [`\u774E`].string() // U+774E <cjk>
	0xF3: [`\u775C`].string() // U+775C <cjk>
	0xF4: [`\u775F`].string() // U+775F <cjk>
	0xF5: [`\u7762`].string() // U+7762 <cjk>
	0xF6: [`\u777A`].string() // U+777A <cjk>
	0xF7: [`\u7780`].string() // U+7780 <cjk>
	0xF8: [`\u7794`].string() // U+7794 <cjk>
	0xF9: [`\u77AA`].string() // U+77AA <cjk>
	0xFA: [`\u77E0`].string() // U+77E0 <cjk>
	0xFB: [`\u782D`].string() // U+782D <cjk>
	0xFC: utf32_to_str(0x2548E) // U+2548E <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x89 = {
	0x40: [`\u9662`].string() // U+9662 <cjk>
	0x41: [`\u9670`].string() // U+9670 <cjk>
	0x42: [`\u96A0`].string() // U+96A0 <cjk>
	0x43: [`\u97FB`].string() // U+97FB <cjk>
	0x44: [`\u540B`].string() // U+540B <cjk>
	0x45: [`\u53F3`].string() // U+53F3 <cjk>
	0x46: [`\u5B87`].string() // U+5B87 <cjk>
	0x47: [`\u70CF`].string() // U+70CF <cjk>
	0x48: [`\u7FBD`].string() // U+7FBD <cjk>
	0x49: [`\u8FC2`].string() // U+8FC2 <cjk>
	0x4A: [`\u96E8`].string() // U+96E8 <cjk>
	0x4B: [`\u536F`].string() // U+536F <cjk>
	0x4C: [`\u9D5C`].string() // U+9D5C <cjk>
	0x4D: [`\u7ABA`].string() // U+7ABA <cjk>
	0x4E: [`\u4E11`].string() // U+4E11 <cjk>
	0x4F: [`\u7893`].string() // U+7893 <cjk>
	0x50: [`\u81FC`].string() // U+81FC <cjk>
	0x51: [`\u6E26`].string() // U+6E26 <cjk>
	0x52: [`\u5618`].string() // U+5618 <cjk>
	0x53: [`\u5504`].string() // U+5504 <cjk>
	0x54: [`\u6B1D`].string() // U+6B1D <cjk>
	0x55: [`\u851A`].string() // U+851A <cjk>
	0x56: [`\u9C3B`].string() // U+9C3B <cjk>
	0x57: [`\u59E5`].string() // U+59E5 <cjk>
	0x58: [`\u53A9`].string() // U+53A9 <cjk>
	0x59: [`\u6D66`].string() // U+6D66 <cjk>
	0x5A: [`\u74DC`].string() // U+74DC <cjk>
	0x5B: [`\u958F`].string() // U+958F <cjk>
	0x5C: [`\u5642`].string() // U+5642 <cjk>
	0x5D: [`\u4E91`].string() // U+4E91 <cjk>
	0x5E: [`\u904B`].string() // U+904B <cjk>
	0x5F: [`\u96F2`].string() // U+96F2 <cjk>
	0x60: [`\u834F`].string() // U+834F <cjk>
	0x61: [`\u990C`].string() // U+990C <cjk>
	0x62: [`\u53E1`].string() // U+53E1 <cjk>
	0x63: [`\u55B6`].string() // U+55B6 <cjk>
	0x64: [`\u5B30`].string() // U+5B30 <cjk>
	0x65: [`\u5F71`].string() // U+5F71 <cjk>
	0x66: [`\u6620`].string() // U+6620 <cjk>
	0x67: [`\u66F3`].string() // U+66F3 <cjk>
	0x68: [`\u6804`].string() // U+6804 <cjk>
	0x69: [`\u6C38`].string() // U+6C38 <cjk>
	0x6A: [`\u6CF3`].string() // U+6CF3 <cjk>
	0x6B: [`\u6D29`].string() // U+6D29 <cjk>
	0x6C: [`\u745B`].string() // U+745B <cjk>
	0x6D: [`\u76C8`].string() // U+76C8 <cjk>
	0x6E: [`\u7A4E`].string() // U+7A4E <cjk>
	0x6F: [`\u9834`].string() // U+9834 <cjk>
	0x70: [`\u82F1`].string() // U+82F1 <cjk>
	0x71: [`\u885B`].string() // U+885B <cjk>
	0x72: [`\u8A60`].string() // U+8A60 <cjk>
	0x73: [`\u92ED`].string() // U+92ED <cjk>
	0x74: [`\u6DB2`].string() // U+6DB2 <cjk>
	0x75: [`\u75AB`].string() // U+75AB <cjk>
	0x76: [`\u76CA`].string() // U+76CA <cjk>
	0x77: [`\u99C5`].string() // U+99C5 <cjk>
	0x78: [`\u60A6`].string() // U+60A6 <cjk>
	0x79: [`\u8B01`].string() // U+8B01 <cjk>
	0x7A: [`\u8D8A`].string() // U+8D8A <cjk>
	0x7B: [`\u95B2`].string() // U+95B2 <cjk>
	0x7C: [`\u698E`].string() // U+698E <cjk>
	0x7D: [`\u53AD`].string() // U+53AD <cjk>
	0x7E: [`\u5186`].string() // U+5186 <cjk>
	0x80: [`\u5712`].string() // U+5712 <cjk>
	0x81: [`\u5830`].string() // U+5830 <cjk>
	0x82: [`\u5944`].string() // U+5944 <cjk>
	0x83: [`\u5BB4`].string() // U+5BB4 <cjk>
	0x84: [`\u5EF6`].string() // U+5EF6 <cjk>
	0x85: [`\u6028`].string() // U+6028 <cjk>
	0x86: [`\u63A9`].string() // U+63A9 <cjk>
	0x87: [`\u63F4`].string() // U+63F4 <cjk>
	0x88: [`\u6CBF`].string() // U+6CBF <cjk>
	0x89: [`\u6F14`].string() // U+6F14 <cjk>
	0x8A: [`\u708E`].string() // U+708E <cjk>
	0x8B: [`\u7114`].string() // U+7114 <cjk>
	0x8C: [`\u7159`].string() // U+7159 <cjk>
	0x8D: [`\u71D5`].string() // U+71D5 <cjk>
	0x8E: [`\u733F`].string() // U+733F <cjk>
	0x8F: [`\u7E01`].string() // U+7E01 <cjk>
	0x90: [`\u8276`].string() // U+8276 <cjk>
	0x91: [`\u82D1`].string() // U+82D1 <cjk>
	0x92: [`\u8597`].string() // U+8597 <cjk>
	0x93: [`\u9060`].string() // U+9060 <cjk>
	0x94: [`\u925B`].string() // U+925B <cjk>
	0x95: [`\u9D1B`].string() // U+9D1B <cjk>
	0x96: [`\u5869`].string() // U+5869 <cjk>
	0x97: [`\u65BC`].string() // U+65BC <cjk>
	0x98: [`\u6C5A`].string() // U+6C5A <cjk>
	0x99: [`\u7525`].string() // U+7525 <cjk>
	0x9A: [`\u51F9`].string() // U+51F9 <cjk>
	0x9B: [`\u592E`].string() // U+592E <cjk>
	0x9C: [`\u5965`].string() // U+5965 <cjk>
	0x9D: [`\u5F80`].string() // U+5F80 <cjk>
	0x9E: [`\u5FDC`].string() // U+5FDC <cjk>
	0x9F: [`\u62BC`].string() // U+62BC <cjk>
	0xA0: [`\u65FA`].string() // U+65FA <cjk>
	0xA1: [`\u6A2A`].string() // U+6A2A <cjk>
	0xA2: [`\u6B27`].string() // U+6B27 <cjk>
	0xA3: [`\u6BB4`].string() // U+6BB4 <cjk>
	0xA4: [`\u738B`].string() // U+738B <cjk>
	0xA5: [`\u7FC1`].string() // U+7FC1 <cjk>
	0xA6: [`\u8956`].string() // U+8956 <cjk>
	0xA7: [`\u9D2C`].string() // U+9D2C <cjk>
	0xA8: [`\u9D0E`].string() // U+9D0E <cjk>
	0xA9: [`\u9EC4`].string() // U+9EC4 <cjk>
	0xAA: [`\u5CA1`].string() // U+5CA1 <cjk>
	0xAB: [`\u6C96`].string() // U+6C96 <cjk>
	0xAC: [`\u837B`].string() // U+837B <cjk>
	0xAD: [`\u5104`].string() // U+5104 <cjk>
	0xAE: [`\u5C4B`].string() // U+5C4B <cjk>
	0xAF: [`\u61B6`].string() // U+61B6 <cjk>
	0xB0: [`\u81C6`].string() // U+81C6 <cjk>
	0xB1: [`\u6876`].string() // U+6876 <cjk>
	0xB2: [`\u7261`].string() // U+7261 <cjk>
	0xB3: [`\u4E59`].string() // U+4E59 <cjk>
	0xB4: [`\u4FFA`].string() // U+4FFA <cjk>
	0xB5: [`\u5378`].string() // U+5378 <cjk>
	0xB6: [`\u6069`].string() // U+6069 <cjk>
	0xB7: [`\u6E29`].string() // U+6E29 <cjk>
	0xB8: [`\u7A4F`].string() // U+7A4F <cjk>
	0xB9: [`\u97F3`].string() // U+97F3 <cjk>
	0xBA: [`\u4E0B`].string() // U+4E0B <cjk>
	0xBB: [`\u5316`].string() // U+5316 <cjk>
	0xBC: [`\u4EEE`].string() // U+4EEE <cjk>
	0xBD: [`\u4F55`].string() // U+4F55 <cjk>
	0xBE: [`\u4F3D`].string() // U+4F3D <cjk>
	0xBF: [`\u4FA1`].string() // U+4FA1 <cjk>
	0xC0: [`\u4F73`].string() // U+4F73 <cjk>
	0xC1: [`\u52A0`].string() // U+52A0 <cjk>
	0xC2: [`\u53EF`].string() // U+53EF <cjk>
	0xC3: [`\u5609`].string() // U+5609 <cjk>
	0xC4: [`\u590F`].string() // U+590F <cjk>
	0xC5: [`\u5AC1`].string() // U+5AC1 <cjk>
	0xC6: [`\u5BB6`].string() // U+5BB6 <cjk>
	0xC7: [`\u5BE1`].string() // U+5BE1 <cjk>
	0xC8: [`\u79D1`].string() // U+79D1 <cjk>
	0xC9: [`\u6687`].string() // U+6687 <cjk>
	0xCA: [`\u679C`].string() // U+679C <cjk>
	0xCB: [`\u67B6`].string() // U+67B6 <cjk>
	0xCC: [`\u6B4C`].string() // U+6B4C <cjk>
	0xCD: [`\u6CB3`].string() // U+6CB3 <cjk>
	0xCE: [`\u706B`].string() // U+706B <cjk>
	0xCF: [`\u73C2`].string() // U+73C2 <cjk>
	0xD0: [`\u798D`].string() // U+798D <cjk>
	0xD1: [`\u79BE`].string() // U+79BE <cjk>
	0xD2: [`\u7A3C`].string() // U+7A3C <cjk>
	0xD3: [`\u7B87`].string() // U+7B87 <cjk>
	0xD4: [`\u82B1`].string() // U+82B1 <cjk>
	0xD5: [`\u82DB`].string() // U+82DB <cjk>
	0xD6: [`\u8304`].string() // U+8304 <cjk>
	0xD7: [`\u8377`].string() // U+8377 <cjk>
	0xD8: [`\u83EF`].string() // U+83EF <cjk>
	0xD9: [`\u83D3`].string() // U+83D3 <cjk>
	0xDA: [`\u8766`].string() // U+8766 <cjk>
	0xDB: [`\u8AB2`].string() // U+8AB2 <cjk>
	0xDC: [`\u5629`].string() // U+5629 <cjk>
	0xDD: [`\u8CA8`].string() // U+8CA8 <cjk>
	0xDE: [`\u8FE6`].string() // U+8FE6 <cjk>
	0xDF: [`\u904E`].string() // U+904E <cjk>
	0xE0: [`\u971E`].string() // U+971E <cjk>
	0xE1: [`\u868A`].string() // U+868A <cjk>
	0xE2: [`\u4FC4`].string() // U+4FC4 <cjk>
	0xE3: [`\u5CE8`].string() // U+5CE8 <cjk>
	0xE4: [`\u6211`].string() // U+6211 <cjk>
	0xE5: [`\u7259`].string() // U+7259 <cjk>
	0xE6: [`\u753B`].string() // U+753B <cjk>
	0xE7: [`\u81E5`].string() // U+81E5 <cjk>
	0xE8: [`\u82BD`].string() // U+82BD <cjk>
	0xE9: [`\u86FE`].string() // U+86FE <cjk>
	0xEA: [`\u8CC0`].string() // U+8CC0 <cjk>
	0xEB: [`\u96C5`].string() // U+96C5 <cjk>
	0xEC: [`\u9913`].string() // U+9913 <cjk>
	0xED: [`\u99D5`].string() // U+99D5 <cjk>
	0xEE: [`\u4ECB`].string() // U+4ECB <cjk>
	0xEF: [`\u4F1A`].string() // U+4F1A <cjk>
	0xF0: [`\u89E3`].string() // U+89E3 <cjk>
	0xF1: [`\u56DE`].string() // U+56DE <cjk>
	0xF2: [`\u584A`].string() // U+584A <cjk>
	0xF3: [`\u58CA`].string() // U+58CA <cjk>
	0xF4: [`\u5EFB`].string() // U+5EFB <cjk>
	0xF5: [`\u5FEB`].string() // U+5FEB <cjk>
	0xF6: [`\u602A`].string() // U+602A <cjk>
	0xF7: [`\u6094`].string() // U+6094 <cjk>
	0xF8: [`\u6062`].string() // U+6062 <cjk>
	0xF9: [`\u61D0`].string() // U+61D0 <cjk>
	0xFA: [`\u6212`].string() // U+6212 <cjk>
	0xFB: [`\u62D0`].string() // U+62D0 <cjk>
	0xFC: [`\u6539`].string() // U+6539 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x9c = {
	0x40: [`\u5ED6`].string() // U+5ED6 <cjk>
	0x41: [`\u5EE3`].string() // U+5EE3 <cjk>
	0x42: [`\u5EDD`].string() // U+5EDD <cjk>
	0x43: [`\u5EDA`].string() // U+5EDA <cjk>
	0x44: [`\u5EDB`].string() // U+5EDB <cjk>
	0x45: [`\u5EE2`].string() // U+5EE2 <cjk>
	0x46: [`\u5EE1`].string() // U+5EE1 <cjk>
	0x47: [`\u5EE8`].string() // U+5EE8 <cjk>
	0x48: [`\u5EE9`].string() // U+5EE9 <cjk>
	0x49: [`\u5EEC`].string() // U+5EEC <cjk>
	0x4A: [`\u5EF1`].string() // U+5EF1 <cjk>
	0x4B: [`\u5EF3`].string() // U+5EF3 <cjk>
	0x4C: [`\u5EF0`].string() // U+5EF0 <cjk>
	0x4D: [`\u5EF4`].string() // U+5EF4 <cjk>
	0x4E: [`\u5EF8`].string() // U+5EF8 <cjk>
	0x4F: [`\u5EFE`].string() // U+5EFE <cjk>
	0x50: [`\u5F03`].string() // U+5F03 <cjk>
	0x51: [`\u5F09`].string() // U+5F09 <cjk>
	0x52: [`\u5F5D`].string() // U+5F5D <cjk>
	0x53: [`\u5F5C`].string() // U+5F5C <cjk>
	0x54: [`\u5F0B`].string() // U+5F0B <cjk>
	0x55: [`\u5F11`].string() // U+5F11 <cjk>
	0x56: [`\u5F16`].string() // U+5F16 <cjk>
	0x57: [`\u5F29`].string() // U+5F29 <cjk>
	0x58: [`\u5F2D`].string() // U+5F2D <cjk>
	0x59: [`\u5F38`].string() // U+5F38 <cjk>
	0x5A: [`\u5F41`].string() // U+5F41 <cjk>
	0x5B: [`\u5F48`].string() // U+5F48 <cjk>
	0x5C: [`\u5F4C`].string() // U+5F4C <cjk>
	0x5D: [`\u5F4E`].string() // U+5F4E <cjk>
	0x5E: [`\u5F2F`].string() // U+5F2F <cjk>
	0x5F: [`\u5F51`].string() // U+5F51 <cjk>
	0x60: [`\u5F56`].string() // U+5F56 <cjk>
	0x61: [`\u5F57`].string() // U+5F57 <cjk>
	0x62: [`\u5F59`].string() // U+5F59 <cjk>
	0x63: [`\u5F61`].string() // U+5F61 <cjk>
	0x64: [`\u5F6D`].string() // U+5F6D <cjk>
	0x65: [`\u5F73`].string() // U+5F73 <cjk>
	0x66: [`\u5F77`].string() // U+5F77 <cjk>
	0x67: [`\u5F83`].string() // U+5F83 <cjk>
	0x68: [`\u5F82`].string() // U+5F82 <cjk>
	0x69: [`\u5F7F`].string() // U+5F7F <cjk>
	0x6A: [`\u5F8A`].string() // U+5F8A <cjk>
	0x6B: [`\u5F88`].string() // U+5F88 <cjk>
	0x6C: [`\u5F91`].string() // U+5F91 <cjk>
	0x6D: [`\u5F87`].string() // U+5F87 <cjk>
	0x6E: [`\u5F9E`].string() // U+5F9E <cjk>
	0x6F: [`\u5F99`].string() // U+5F99 <cjk>
	0x70: [`\u5F98`].string() // U+5F98 <cjk>
	0x71: [`\u5FA0`].string() // U+5FA0 <cjk>
	0x72: [`\u5FA8`].string() // U+5FA8 <cjk>
	0x73: [`\u5FAD`].string() // U+5FAD <cjk>
	0x74: [`\u5FBC`].string() // U+5FBC <cjk>
	0x75: [`\u5FD6`].string() // U+5FD6 <cjk>
	0x76: [`\u5FFB`].string() // U+5FFB <cjk>
	0x77: [`\u5FE4`].string() // U+5FE4 <cjk>
	0x78: [`\u5FF8`].string() // U+5FF8 <cjk>
	0x79: [`\u5FF1`].string() // U+5FF1 <cjk>
	0x7A: [`\u5FDD`].string() // U+5FDD <cjk>
	0x7B: [`\u60B3`].string() // U+60B3 <cjk>
	0x7C: [`\u5FFF`].string() // U+5FFF <cjk>
	0x7D: [`\u6021`].string() // U+6021 <cjk>
	0x7E: [`\u6060`].string() // U+6060 <cjk>
	0x80: [`\u6019`].string() // U+6019 <cjk>
	0x81: [`\u6010`].string() // U+6010 <cjk>
	0x82: [`\u6029`].string() // U+6029 <cjk>
	0x83: [`\u600E`].string() // U+600E <cjk>
	0x84: [`\u6031`].string() // U+6031 <cjk>
	0x85: [`\u601B`].string() // U+601B <cjk>
	0x86: [`\u6015`].string() // U+6015 <cjk>
	0x87: [`\u602B`].string() // U+602B <cjk>
	0x88: [`\u6026`].string() // U+6026 <cjk>
	0x89: [`\u600F`].string() // U+600F <cjk>
	0x8A: [`\u603A`].string() // U+603A <cjk>
	0x8B: [`\u605A`].string() // U+605A <cjk>
	0x8C: [`\u6041`].string() // U+6041 <cjk>
	0x8D: [`\u606A`].string() // U+606A <cjk>
	0x8E: [`\u6077`].string() // U+6077 <cjk>
	0x8F: [`\u605F`].string() // U+605F <cjk>
	0x90: [`\u604A`].string() // U+604A <cjk>
	0x91: [`\u6046`].string() // U+6046 <cjk>
	0x92: [`\u604D`].string() // U+604D <cjk>
	0x93: [`\u6063`].string() // U+6063 <cjk>
	0x94: [`\u6043`].string() // U+6043 <cjk>
	0x95: [`\u6064`].string() // U+6064 <cjk>
	0x96: [`\u6042`].string() // U+6042 <cjk>
	0x97: [`\u606C`].string() // U+606C <cjk>
	0x98: [`\u606B`].string() // U+606B <cjk>
	0x99: [`\u6059`].string() // U+6059 <cjk>
	0x9A: [`\u6081`].string() // U+6081 <cjk>
	0x9B: [`\u608D`].string() // U+608D <cjk>
	0x9C: [`\u60E7`].string() // U+60E7 <cjk>
	0x9D: [`\u6083`].string() // U+6083 <cjk>
	0x9E: [`\u609A`].string() // U+609A <cjk>
	0x9F: [`\u6084`].string() // U+6084 <cjk>
	0xA0: [`\u609B`].string() // U+609B <cjk>
	0xA1: [`\u6096`].string() // U+6096 <cjk>
	0xA2: [`\u6097`].string() // U+6097 <cjk>
	0xA3: [`\u6092`].string() // U+6092 <cjk>
	0xA4: [`\u60A7`].string() // U+60A7 <cjk>
	0xA5: [`\u608B`].string() // U+608B <cjk>
	0xA6: [`\u60E1`].string() // U+60E1 <cjk>
	0xA7: [`\u60B8`].string() // U+60B8 <cjk>
	0xA8: [`\u60E0`].string() // U+60E0 <cjk>
	0xA9: [`\u60D3`].string() // U+60D3 <cjk>
	0xAA: [`\u60B4`].string() // U+60B4 <cjk>
	0xAB: [`\u5FF0`].string() // U+5FF0 <cjk>
	0xAC: [`\u60BD`].string() // U+60BD <cjk>
	0xAD: [`\u60C6`].string() // U+60C6 <cjk>
	0xAE: [`\u60B5`].string() // U+60B5 <cjk>
	0xAF: [`\u60D8`].string() // U+60D8 <cjk>
	0xB0: [`\u614D`].string() // U+614D <cjk>
	0xB1: [`\u6115`].string() // U+6115 <cjk>
	0xB2: [`\u6106`].string() // U+6106 <cjk>
	0xB3: [`\u60F6`].string() // U+60F6 <cjk>
	0xB4: [`\u60F7`].string() // U+60F7 <cjk>
	0xB5: [`\u6100`].string() // U+6100 <cjk>
	0xB6: [`\u60F4`].string() // U+60F4 <cjk>
	0xB7: [`\u60FA`].string() // U+60FA <cjk>
	0xB8: [`\u6103`].string() // U+6103 <cjk>
	0xB9: [`\u6121`].string() // U+6121 <cjk>
	0xBA: [`\u60FB`].string() // U+60FB <cjk>
	0xBB: [`\u60F1`].string() // U+60F1 <cjk>
	0xBC: [`\u610D`].string() // U+610D <cjk>
	0xBD: [`\u610E`].string() // U+610E <cjk>
	0xBE: [`\u6147`].string() // U+6147 <cjk>
	0xBF: [`\u613E`].string() // U+613E <cjk>
	0xC0: [`\u6128`].string() // U+6128 <cjk>
	0xC1: [`\u6127`].string() // U+6127 <cjk>
	0xC2: [`\u614A`].string() // U+614A <cjk>
	0xC3: [`\u613F`].string() // U+613F <cjk>
	0xC4: [`\u613C`].string() // U+613C <cjk>
	0xC5: [`\u612C`].string() // U+612C <cjk>
	0xC6: [`\u6134`].string() // U+6134 <cjk>
	0xC7: [`\u613D`].string() // U+613D <cjk>
	0xC8: [`\u6142`].string() // U+6142 <cjk>
	0xC9: [`\u6144`].string() // U+6144 <cjk>
	0xCA: [`\u6173`].string() // U+6173 <cjk>
	0xCB: [`\u6177`].string() // U+6177 <cjk>
	0xCC: [`\u6158`].string() // U+6158 <cjk>
	0xCD: [`\u6159`].string() // U+6159 <cjk>
	0xCE: [`\u615A`].string() // U+615A <cjk>
	0xCF: [`\u616B`].string() // U+616B <cjk>
	0xD0: [`\u6174`].string() // U+6174 <cjk>
	0xD1: [`\u616F`].string() // U+616F <cjk>
	0xD2: [`\u6165`].string() // U+6165 <cjk>
	0xD3: [`\u6171`].string() // U+6171 <cjk>
	0xD4: [`\u615F`].string() // U+615F <cjk>
	0xD5: [`\u615D`].string() // U+615D <cjk>
	0xD6: [`\u6153`].string() // U+6153 <cjk>
	0xD7: [`\u6175`].string() // U+6175 <cjk>
	0xD8: [`\u6199`].string() // U+6199 <cjk>
	0xD9: [`\u6196`].string() // U+6196 <cjk>
	0xDA: [`\u6187`].string() // U+6187 <cjk>
	0xDB: [`\u61AC`].string() // U+61AC <cjk>
	0xDC: [`\u6194`].string() // U+6194 <cjk>
	0xDD: [`\u619A`].string() // U+619A <cjk>
	0xDE: [`\u618A`].string() // U+618A <cjk>
	0xDF: [`\u6191`].string() // U+6191 <cjk>
	0xE0: [`\u61AB`].string() // U+61AB <cjk>
	0xE1: [`\u61AE`].string() // U+61AE <cjk>
	0xE2: [`\u61CC`].string() // U+61CC <cjk>
	0xE3: [`\u61CA`].string() // U+61CA <cjk>
	0xE4: [`\u61C9`].string() // U+61C9 <cjk>
	0xE5: [`\u61F7`].string() // U+61F7 <cjk>
	0xE6: [`\u61C8`].string() // U+61C8 <cjk>
	0xE7: [`\u61C3`].string() // U+61C3 <cjk>
	0xE8: [`\u61C6`].string() // U+61C6 <cjk>
	0xE9: [`\u61BA`].string() // U+61BA <cjk>
	0xEA: [`\u61CB`].string() // U+61CB <cjk>
	0xEB: [`\u7F79`].string() // U+7F79 <cjk>
	0xEC: [`\u61CD`].string() // U+61CD <cjk>
	0xED: [`\u61E6`].string() // U+61E6 <cjk>
	0xEE: [`\u61E3`].string() // U+61E3 <cjk>
	0xEF: [`\u61F6`].string() // U+61F6 <cjk>
	0xF0: [`\u61FA`].string() // U+61FA <cjk>
	0xF1: [`\u61F4`].string() // U+61F4 <cjk>
	0xF2: [`\u61FF`].string() // U+61FF <cjk>
	0xF3: [`\u61FD`].string() // U+61FD <cjk>
	0xF4: [`\u61FC`].string() // U+61FC <cjk>
	0xF5: [`\u61FE`].string() // U+61FE <cjk>
	0xF6: [`\u6200`].string() // U+6200 <cjk>
	0xF7: [`\u6208`].string() // U+6208 <cjk>
	0xF8: [`\u6209`].string() // U+6209 <cjk>
	0xF9: [`\u620D`].string() // U+620D <cjk>
	0xFA: [`\u620C`].string() // U+620C <cjk>
	0xFB: [`\u6214`].string() // U+6214 <cjk>
	0xFC: [`\u621B`].string() // U+621B <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xe6 = {
	0x40: [`\u8966`].string() // U+8966 <cjk>
	0x41: [`\u8964`].string() // U+8964 <cjk>
	0x42: [`\u896D`].string() // U+896D <cjk>
	0x43: [`\u896A`].string() // U+896A <cjk>
	0x44: [`\u896F`].string() // U+896F <cjk>
	0x45: [`\u8974`].string() // U+8974 <cjk>
	0x46: [`\u8977`].string() // U+8977 <cjk>
	0x47: [`\u897E`].string() // U+897E <cjk>
	0x48: [`\u8983`].string() // U+8983 <cjk>
	0x49: [`\u8988`].string() // U+8988 <cjk>
	0x4A: [`\u898A`].string() // U+898A <cjk>
	0x4B: [`\u8993`].string() // U+8993 <cjk>
	0x4C: [`\u8998`].string() // U+8998 <cjk>
	0x4D: [`\u89A1`].string() // U+89A1 <cjk>
	0x4E: [`\u89A9`].string() // U+89A9 <cjk>
	0x4F: [`\u89A6`].string() // U+89A6 <cjk>
	0x50: [`\u89AC`].string() // U+89AC <cjk>
	0x51: [`\u89AF`].string() // U+89AF <cjk>
	0x52: [`\u89B2`].string() // U+89B2 <cjk>
	0x53: [`\u89BA`].string() // U+89BA <cjk>
	0x54: [`\u89BD`].string() // U+89BD <cjk>
	0x55: [`\u89BF`].string() // U+89BF <cjk>
	0x56: [`\u89C0`].string() // U+89C0 <cjk>
	0x57: [`\u89DA`].string() // U+89DA <cjk>
	0x58: [`\u89DC`].string() // U+89DC <cjk>
	0x59: [`\u89DD`].string() // U+89DD <cjk>
	0x5A: [`\u89E7`].string() // U+89E7 <cjk>
	0x5B: [`\u89F4`].string() // U+89F4 <cjk>
	0x5C: [`\u89F8`].string() // U+89F8 <cjk>
	0x5D: [`\u8A03`].string() // U+8A03 <cjk>
	0x5E: [`\u8A16`].string() // U+8A16 <cjk>
	0x5F: [`\u8A10`].string() // U+8A10 <cjk>
	0x60: [`\u8A0C`].string() // U+8A0C <cjk>
	0x61: [`\u8A1B`].string() // U+8A1B <cjk>
	0x62: [`\u8A1D`].string() // U+8A1D <cjk>
	0x63: [`\u8A25`].string() // U+8A25 <cjk>
	0x64: [`\u8A36`].string() // U+8A36 <cjk>
	0x65: [`\u8A41`].string() // U+8A41 <cjk>
	0x66: [`\u8A5B`].string() // U+8A5B <cjk>
	0x67: [`\u8A52`].string() // U+8A52 <cjk>
	0x68: [`\u8A46`].string() // U+8A46 <cjk>
	0x69: [`\u8A48`].string() // U+8A48 <cjk>
	0x6A: [`\u8A7C`].string() // U+8A7C <cjk>
	0x6B: [`\u8A6D`].string() // U+8A6D <cjk>
	0x6C: [`\u8A6C`].string() // U+8A6C <cjk>
	0x6D: [`\u8A62`].string() // U+8A62 <cjk>
	0x6E: [`\u8A85`].string() // U+8A85 <cjk>
	0x6F: [`\u8A82`].string() // U+8A82 <cjk>
	0x70: [`\u8A84`].string() // U+8A84 <cjk>
	0x71: [`\u8AA8`].string() // U+8AA8 <cjk>
	0x72: [`\u8AA1`].string() // U+8AA1 <cjk>
	0x73: [`\u8A91`].string() // U+8A91 <cjk>
	0x74: [`\u8AA5`].string() // U+8AA5 <cjk>
	0x75: [`\u8AA6`].string() // U+8AA6 <cjk>
	0x76: [`\u8A9A`].string() // U+8A9A <cjk>
	0x77: [`\u8AA3`].string() // U+8AA3 <cjk>
	0x78: [`\u8AC4`].string() // U+8AC4 <cjk>
	0x79: [`\u8ACD`].string() // U+8ACD <cjk>
	0x7A: [`\u8AC2`].string() // U+8AC2 <cjk>
	0x7B: [`\u8ADA`].string() // U+8ADA <cjk>
	0x7C: [`\u8AEB`].string() // U+8AEB <cjk>
	0x7D: [`\u8AF3`].string() // U+8AF3 <cjk>
	0x7E: [`\u8AE7`].string() // U+8AE7 <cjk>
	0x80: [`\u8AE4`].string() // U+8AE4 <cjk>
	0x81: [`\u8AF1`].string() // U+8AF1 <cjk>
	0x82: [`\u8B14`].string() // U+8B14 <cjk>
	0x83: [`\u8AE0`].string() // U+8AE0 <cjk>
	0x84: [`\u8AE2`].string() // U+8AE2 <cjk>
	0x85: [`\u8AF7`].string() // U+8AF7 <cjk>
	0x86: [`\u8ADE`].string() // U+8ADE <cjk>
	0x87: [`\u8ADB`].string() // U+8ADB <cjk>
	0x88: [`\u8B0C`].string() // U+8B0C <cjk>
	0x89: [`\u8B07`].string() // U+8B07 <cjk>
	0x8A: [`\u8B1A`].string() // U+8B1A <cjk>
	0x8B: [`\u8AE1`].string() // U+8AE1 <cjk>
	0x8C: [`\u8B16`].string() // U+8B16 <cjk>
	0x8D: [`\u8B10`].string() // U+8B10 <cjk>
	0x8E: [`\u8B17`].string() // U+8B17 <cjk>
	0x8F: [`\u8B20`].string() // U+8B20 <cjk>
	0x90: [`\u8B33`].string() // U+8B33 <cjk>
	0x91: [`\u97AB`].string() // U+97AB <cjk>
	0x92: [`\u8B26`].string() // U+8B26 <cjk>
	0x93: [`\u8B2B`].string() // U+8B2B <cjk>
	0x94: [`\u8B3E`].string() // U+8B3E <cjk>
	0x95: [`\u8B28`].string() // U+8B28 <cjk>
	0x96: [`\u8B41`].string() // U+8B41 <cjk>
	0x97: [`\u8B4C`].string() // U+8B4C <cjk>
	0x98: [`\u8B4F`].string() // U+8B4F <cjk>
	0x99: [`\u8B4E`].string() // U+8B4E <cjk>
	0x9A: [`\u8B49`].string() // U+8B49 <cjk>
	0x9B: [`\u8B56`].string() // U+8B56 <cjk>
	0x9C: [`\u8B5B`].string() // U+8B5B <cjk>
	0x9D: [`\u8B5A`].string() // U+8B5A <cjk>
	0x9E: [`\u8B6B`].string() // U+8B6B <cjk>
	0x9F: [`\u8B5F`].string() // U+8B5F <cjk>
	0xA0: [`\u8B6C`].string() // U+8B6C <cjk>
	0xA1: [`\u8B6F`].string() // U+8B6F <cjk>
	0xA2: [`\u8B74`].string() // U+8B74 <cjk>
	0xA3: [`\u8B7D`].string() // U+8B7D <cjk>
	0xA4: [`\u8B80`].string() // U+8B80 <cjk>
	0xA5: [`\u8B8C`].string() // U+8B8C <cjk>
	0xA6: [`\u8B8E`].string() // U+8B8E <cjk>
	0xA7: [`\u8B92`].string() // U+8B92 <cjk>
	0xA8: [`\u8B93`].string() // U+8B93 <cjk>
	0xA9: [`\u8B96`].string() // U+8B96 <cjk>
	0xAA: [`\u8B99`].string() // U+8B99 <cjk>
	0xAB: [`\u8B9A`].string() // U+8B9A <cjk>
	0xAC: [`\u8C3A`].string() // U+8C3A <cjk>
	0xAD: [`\u8C41`].string() // U+8C41 <cjk>
	0xAE: [`\u8C3F`].string() // U+8C3F <cjk>
	0xAF: [`\u8C48`].string() // U+8C48 <cjk>
	0xB0: [`\u8C4C`].string() // U+8C4C <cjk>
	0xB1: [`\u8C4E`].string() // U+8C4E <cjk>
	0xB2: [`\u8C50`].string() // U+8C50 <cjk>
	0xB3: [`\u8C55`].string() // U+8C55 <cjk>
	0xB4: [`\u8C62`].string() // U+8C62 <cjk>
	0xB5: [`\u8C6C`].string() // U+8C6C <cjk>
	0xB6: [`\u8C78`].string() // U+8C78 <cjk>
	0xB7: [`\u8C7A`].string() // U+8C7A <cjk>
	0xB8: [`\u8C82`].string() // U+8C82 <cjk>
	0xB9: [`\u8C89`].string() // U+8C89 <cjk>
	0xBA: [`\u8C85`].string() // U+8C85 <cjk>
	0xBB: [`\u8C8A`].string() // U+8C8A <cjk>
	0xBC: [`\u8C8D`].string() // U+8C8D <cjk>
	0xBD: [`\u8C8E`].string() // U+8C8E <cjk>
	0xBE: [`\u8C94`].string() // U+8C94 <cjk>
	0xBF: [`\u8C7C`].string() // U+8C7C <cjk>
	0xC0: [`\u8C98`].string() // U+8C98 <cjk>
	0xC1: [`\u621D`].string() // U+621D <cjk>
	0xC2: [`\u8CAD`].string() // U+8CAD <cjk>
	0xC3: [`\u8CAA`].string() // U+8CAA <cjk>
	0xC4: [`\u8CBD`].string() // U+8CBD <cjk>
	0xC5: [`\u8CB2`].string() // U+8CB2 <cjk>
	0xC6: [`\u8CB3`].string() // U+8CB3 <cjk>
	0xC7: [`\u8CAE`].string() // U+8CAE <cjk>
	0xC8: [`\u8CB6`].string() // U+8CB6 <cjk>
	0xC9: [`\u8CC8`].string() // U+8CC8 <cjk>
	0xCA: [`\u8CC1`].string() // U+8CC1 <cjk>
	0xCB: [`\u8CE4`].string() // U+8CE4 <cjk>
	0xCC: [`\u8CE3`].string() // U+8CE3 <cjk>
	0xCD: [`\u8CDA`].string() // U+8CDA <cjk>
	0xCE: [`\u8CFD`].string() // U+8CFD <cjk>
	0xCF: [`\u8CFA`].string() // U+8CFA <cjk>
	0xD0: [`\u8CFB`].string() // U+8CFB <cjk>
	0xD1: [`\u8D04`].string() // U+8D04 <cjk>
	0xD2: [`\u8D05`].string() // U+8D05 <cjk>
	0xD3: [`\u8D0A`].string() // U+8D0A <cjk>
	0xD4: [`\u8D07`].string() // U+8D07 <cjk>
	0xD5: [`\u8D0F`].string() // U+8D0F <cjk>
	0xD6: [`\u8D0D`].string() // U+8D0D <cjk>
	0xD7: [`\u8D10`].string() // U+8D10 <cjk>
	0xD8: [`\u9F4E`].string() // U+9F4E <cjk>
	0xD9: [`\u8D13`].string() // U+8D13 <cjk>
	0xDA: [`\u8CCD`].string() // U+8CCD <cjk>
	0xDB: [`\u8D14`].string() // U+8D14 <cjk>
	0xDC: [`\u8D16`].string() // U+8D16 <cjk>
	0xDD: [`\u8D67`].string() // U+8D67 <cjk>
	0xDE: [`\u8D6D`].string() // U+8D6D <cjk>
	0xDF: [`\u8D71`].string() // U+8D71 <cjk>
	0xE0: [`\u8D73`].string() // U+8D73 <cjk>
	0xE1: [`\u8D81`].string() // U+8D81 <cjk>
	0xE2: [`\u8D99`].string() // U+8D99 <cjk>
	0xE3: [`\u8DC2`].string() // U+8DC2 <cjk>
	0xE4: [`\u8DBE`].string() // U+8DBE <cjk>
	0xE5: [`\u8DBA`].string() // U+8DBA <cjk>
	0xE6: [`\u8DCF`].string() // U+8DCF <cjk>
	0xE7: [`\u8DDA`].string() // U+8DDA <cjk>
	0xE8: [`\u8DD6`].string() // U+8DD6 <cjk>
	0xE9: [`\u8DCC`].string() // U+8DCC <cjk>
	0xEA: [`\u8DDB`].string() // U+8DDB <cjk>
	0xEB: [`\u8DCB`].string() // U+8DCB <cjk>
	0xEC: [`\u8DEA`].string() // U+8DEA <cjk>
	0xED: [`\u8DEB`].string() // U+8DEB <cjk>
	0xEE: [`\u8DDF`].string() // U+8DDF <cjk>
	0xEF: [`\u8DE3`].string() // U+8DE3 <cjk>
	0xF0: [`\u8DFC`].string() // U+8DFC <cjk>
	0xF1: [`\u8E08`].string() // U+8E08 <cjk>
	0xF2: [`\u8E09`].string() // U+8E09 <cjk>
	0xF3: [`\u8DFF`].string() // U+8DFF <cjk>
	0xF4: [`\u8E1D`].string() // U+8E1D <cjk>
	0xF5: [`\u8E1E`].string() // U+8E1E <cjk>
	0xF6: [`\u8E10`].string() // U+8E10 <cjk>
	0xF7: [`\u8E1F`].string() // U+8E1F <cjk>
	0xF8: [`\u8E42`].string() // U+8E42 <cjk>
	0xF9: [`\u8E35`].string() // U+8E35 <cjk>
	0xFA: [`\u8E30`].string() // U+8E30 <cjk>
	0xFB: [`\u8E34`].string() // U+8E34 <cjk>
	0xFC: [`\u8E4A`].string() // U+8E4A <cjk>
}

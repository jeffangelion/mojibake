module mojibake

const jis_x_0213_doublebyte_0x8e = {
	0x40: [`\u5BDF`].string() // U+5BDF <cjk>
	0x41: [`\u62F6`].string() // U+62F6 <cjk>
	0x42: [`\u64AE`].string() // U+64AE <cjk>
	0x43: [`\u64E6`].string() // U+64E6 <cjk>
	0x44: [`\u672D`].string() // U+672D <cjk>
	0x45: [`\u6BBA`].string() // U+6BBA <cjk>
	0x46: [`\u85A9`].string() // U+85A9 <cjk>
	0x47: [`\u96D1`].string() // U+96D1 <cjk>
	0x48: [`\u7690`].string() // U+7690 <cjk>
	0x49: [`\u9BD6`].string() // U+9BD6 <cjk>
	0x4A: [`\u634C`].string() // U+634C <cjk>
	0x4B: [`\u9306`].string() // U+9306 <cjk>
	0x4C: [`\u9BAB`].string() // U+9BAB <cjk>
	0x4D: [`\u76BF`].string() // U+76BF <cjk>
	0x4E: [`\u6652`].string() // U+6652 <cjk>
	0x4F: [`\u4E09`].string() // U+4E09 <cjk>
	0x50: [`\u5098`].string() // U+5098 <cjk>
	0x51: [`\u53C2`].string() // U+53C2 <cjk>
	0x52: [`\u5C71`].string() // U+5C71 <cjk>
	0x53: [`\u60E8`].string() // U+60E8 <cjk>
	0x54: [`\u6492`].string() // U+6492 <cjk>
	0x55: [`\u6563`].string() // U+6563 <cjk>
	0x56: [`\u685F`].string() // U+685F <cjk>
	0x57: [`\u71E6`].string() // U+71E6 <cjk>
	0x58: [`\u73CA`].string() // U+73CA <cjk>
	0x59: [`\u7523`].string() // U+7523 <cjk>
	0x5A: [`\u7B97`].string() // U+7B97 <cjk>
	0x5B: [`\u7E82`].string() // U+7E82 <cjk>
	0x5C: [`\u8695`].string() // U+8695 <cjk>
	0x5D: [`\u8B83`].string() // U+8B83 <cjk>
	0x5E: [`\u8CDB`].string() // U+8CDB <cjk>
	0x5F: [`\u9178`].string() // U+9178 <cjk>
	0x60: [`\u9910`].string() // U+9910 <cjk>
	0x61: [`\u65AC`].string() // U+65AC <cjk>
	0x62: [`\u66AB`].string() // U+66AB <cjk>
	0x63: [`\u6B8B`].string() // U+6B8B <cjk>
	0x64: [`\u4ED5`].string() // U+4ED5 <cjk>
	0x65: [`\u4ED4`].string() // U+4ED4 <cjk>
	0x66: [`\u4F3A`].string() // U+4F3A <cjk>
	0x67: [`\u4F7F`].string() // U+4F7F <cjk>
	0x68: [`\u523A`].string() // U+523A <cjk>
	0x69: [`\u53F8`].string() // U+53F8 <cjk>
	0x6A: [`\u53F2`].string() // U+53F2 <cjk>
	0x6B: [`\u55E3`].string() // U+55E3 <cjk>
	0x6C: [`\u56DB`].string() // U+56DB <cjk>
	0x6D: [`\u58EB`].string() // U+58EB <cjk>
	0x6E: [`\u59CB`].string() // U+59CB <cjk>
	0x6F: [`\u59C9`].string() // U+59C9 <cjk>
	0x70: [`\u59FF`].string() // U+59FF <cjk>
	0x71: [`\u5B50`].string() // U+5B50 <cjk>
	0x72: [`\u5C4D`].string() // U+5C4D <cjk>
	0x73: [`\u5E02`].string() // U+5E02 <cjk>
	0x74: [`\u5E2B`].string() // U+5E2B <cjk>
	0x75: [`\u5FD7`].string() // U+5FD7 <cjk>
	0x76: [`\u601D`].string() // U+601D <cjk>
	0x77: [`\u6307`].string() // U+6307 <cjk>
	0x78: [`\u652F`].string() // U+652F <cjk>
	0x79: [`\u5B5C`].string() // U+5B5C <cjk>
	0x7A: [`\u65AF`].string() // U+65AF <cjk>
	0x7B: [`\u65BD`].string() // U+65BD <cjk>
	0x7C: [`\u65E8`].string() // U+65E8 <cjk>
	0x7D: [`\u679D`].string() // U+679D <cjk>
	0x7E: [`\u6B62`].string() // U+6B62 <cjk>
	0x80: [`\u6B7B`].string() // U+6B7B <cjk>
	0x81: [`\u6C0F`].string() // U+6C0F <cjk>
	0x82: [`\u7345`].string() // U+7345 <cjk>
	0x83: [`\u7949`].string() // U+7949 <cjk>
	0x84: [`\u79C1`].string() // U+79C1 <cjk>
	0x85: [`\u7CF8`].string() // U+7CF8 <cjk>
	0x86: [`\u7D19`].string() // U+7D19 <cjk>
	0x87: [`\u7D2B`].string() // U+7D2B <cjk>
	0x88: [`\u80A2`].string() // U+80A2 <cjk>
	0x89: [`\u8102`].string() // U+8102 <cjk>
	0x8A: [`\u81F3`].string() // U+81F3 <cjk>
	0x8B: [`\u8996`].string() // U+8996 <cjk>
	0x8C: [`\u8A5E`].string() // U+8A5E <cjk>
	0x8D: [`\u8A69`].string() // U+8A69 <cjk>
	0x8E: [`\u8A66`].string() // U+8A66 <cjk>
	0x8F: [`\u8A8C`].string() // U+8A8C <cjk>
	0x90: [`\u8AEE`].string() // U+8AEE <cjk>
	0x91: [`\u8CC7`].string() // U+8CC7 <cjk>
	0x92: [`\u8CDC`].string() // U+8CDC <cjk>
	0x93: [`\u96CC`].string() // U+96CC <cjk>
	0x94: [`\u98FC`].string() // U+98FC <cjk>
	0x95: [`\u6B6F`].string() // U+6B6F <cjk>
	0x96: [`\u4E8B`].string() // U+4E8B <cjk>
	0x97: [`\u4F3C`].string() // U+4F3C <cjk>
	0x98: [`\u4F8D`].string() // U+4F8D <cjk>
	0x99: [`\u5150`].string() // U+5150 <cjk>
	0x9A: [`\u5B57`].string() // U+5B57 <cjk>
	0x9B: [`\u5BFA`].string() // U+5BFA <cjk>
	0x9C: [`\u6148`].string() // U+6148 <cjk>
	0x9D: [`\u6301`].string() // U+6301 <cjk>
	0x9E: [`\u6642`].string() // U+6642 <cjk>
	0x9F: [`\u6B21`].string() // U+6B21 <cjk>
	0xA0: [`\u6ECB`].string() // U+6ECB <cjk>
	0xA1: [`\u6CBB`].string() // U+6CBB <cjk>
	0xA2: [`\u723E`].string() // U+723E <cjk>
	0xA3: [`\u74BD`].string() // U+74BD <cjk>
	0xA4: [`\u75D4`].string() // U+75D4 <cjk>
	0xA5: [`\u78C1`].string() // U+78C1 <cjk>
	0xA6: [`\u793A`].string() // U+793A <cjk>
	0xA7: [`\u800C`].string() // U+800C <cjk>
	0xA8: [`\u8033`].string() // U+8033 <cjk>
	0xA9: [`\u81EA`].string() // U+81EA <cjk>
	0xAA: [`\u8494`].string() // U+8494 <cjk>
	0xAB: [`\u8F9E`].string() // U+8F9E <cjk>
	0xAC: [`\u6C50`].string() // U+6C50 <cjk>
	0xAD: [`\u9E7F`].string() // U+9E7F <cjk>
	0xAE: [`\u5F0F`].string() // U+5F0F <cjk>
	0xAF: [`\u8B58`].string() // U+8B58 <cjk>
	0xB0: [`\u9D2B`].string() // U+9D2B <cjk>
	0xB1: [`\u7AFA`].string() // U+7AFA <cjk>
	0xB2: [`\u8EF8`].string() // U+8EF8 <cjk>
	0xB3: [`\u5B8D`].string() // U+5B8D <cjk>
	0xB4: [`\u96EB`].string() // U+96EB <cjk>
	0xB5: [`\u4E03`].string() // U+4E03 <cjk>
	0xB6: [`\u53F1`].string() // U+53F1 <cjk>
	0xB7: [`\u57F7`].string() // U+57F7 <cjk>
	0xB8: [`\u5931`].string() // U+5931 <cjk>
	0xB9: [`\u5AC9`].string() // U+5AC9 <cjk>
	0xBA: [`\u5BA4`].string() // U+5BA4 <cjk>
	0xBB: [`\u6089`].string() // U+6089 <cjk>
	0xBC: [`\u6E7F`].string() // U+6E7F <cjk>
	0xBD: [`\u6F06`].string() // U+6F06 <cjk>
	0xBE: [`\u75BE`].string() // U+75BE <cjk>
	0xBF: [`\u8CEA`].string() // U+8CEA <cjk>
	0xC0: [`\u5B9F`].string() // U+5B9F <cjk>
	0xC1: [`\u8500`].string() // U+8500 <cjk>
	0xC2: [`\u7BE0`].string() // U+7BE0 <cjk>
	0xC3: [`\u5072`].string() // U+5072 <cjk>
	0xC4: [`\u67F4`].string() // U+67F4 <cjk>
	0xC5: [`\u829D`].string() // U+829D <cjk>
	0xC6: [`\u5C61`].string() // U+5C61 <cjk>
	0xC7: [`\u854A`].string() // U+854A <cjk>
	0xC8: [`\u7E1E`].string() // U+7E1E <cjk>
	0xC9: [`\u820E`].string() // U+820E <cjk>
	0xCA: [`\u5199`].string() // U+5199 <cjk>
	0xCB: [`\u5C04`].string() // U+5C04 <cjk>
	0xCC: [`\u6368`].string() // U+6368 <cjk>
	0xCD: [`\u8D66`].string() // U+8D66 <cjk>
	0xCE: [`\u659C`].string() // U+659C <cjk>
	0xCF: [`\u716E`].string() // U+716E <cjk>
	0xD0: [`\u793E`].string() // U+793E <cjk>
	0xD1: [`\u7D17`].string() // U+7D17 <cjk>
	0xD2: [`\u8005`].string() // U+8005 <cjk>
	0xD3: [`\u8B1D`].string() // U+8B1D <cjk>
	0xD4: [`\u8ECA`].string() // U+8ECA <cjk>
	0xD5: [`\u906E`].string() // U+906E <cjk>
	0xD6: [`\u86C7`].string() // U+86C7 <cjk>
	0xD7: [`\u90AA`].string() // U+90AA <cjk>
	0xD8: [`\u501F`].string() // U+501F <cjk>
	0xD9: [`\u52FA`].string() // U+52FA <cjk>
	0xDA: [`\u5C3A`].string() // U+5C3A <cjk>
	0xDB: [`\u6753`].string() // U+6753 <cjk>
	0xDC: [`\u707C`].string() // U+707C <cjk>
	0xDD: [`\u7235`].string() // U+7235 <cjk>
	0xDE: [`\u914C`].string() // U+914C <cjk>
	0xDF: [`\u91C8`].string() // U+91C8 <cjk>
	0xE0: [`\u932B`].string() // U+932B <cjk>
	0xE1: [`\u82E5`].string() // U+82E5 <cjk>
	0xE2: [`\u5BC2`].string() // U+5BC2 <cjk>
	0xE3: [`\u5F31`].string() // U+5F31 <cjk>
	0xE4: [`\u60F9`].string() // U+60F9 <cjk>
	0xE5: [`\u4E3B`].string() // U+4E3B <cjk>
	0xE6: [`\u53D6`].string() // U+53D6 <cjk>
	0xE7: [`\u5B88`].string() // U+5B88 <cjk>
	0xE8: [`\u624B`].string() // U+624B <cjk>
	0xE9: [`\u6731`].string() // U+6731 <cjk>
	0xEA: [`\u6B8A`].string() // U+6B8A <cjk>
	0xEB: [`\u72E9`].string() // U+72E9 <cjk>
	0xEC: [`\u73E0`].string() // U+73E0 <cjk>
	0xED: [`\u7A2E`].string() // U+7A2E <cjk>
	0xEE: [`\u816B`].string() // U+816B <cjk>
	0xEF: [`\u8DA3`].string() // U+8DA3 <cjk>
	0xF0: [`\u9152`].string() // U+9152 <cjk>
	0xF1: [`\u9996`].string() // U+9996 <cjk>
	0xF2: [`\u5112`].string() // U+5112 <cjk>
	0xF3: [`\u53D7`].string() // U+53D7 <cjk>
	0xF4: [`\u546A`].string() // U+546A <cjk>
	0xF5: [`\u5BFF`].string() // U+5BFF <cjk>
	0xF6: [`\u6388`].string() // U+6388 <cjk>
	0xF7: [`\u6A39`].string() // U+6A39 <cjk>
	0xF8: [`\u7DAC`].string() // U+7DAC <cjk>
	0xF9: [`\u9700`].string() // U+9700 <cjk>
	0xFA: [`\u56DA`].string() // U+56DA <cjk>
	0xFB: [`\u53CE`].string() // U+53CE <cjk>
	0xFC: [`\u5468`].string() // U+5468 <cjk>
}

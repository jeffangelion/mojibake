module mojibake

const jis_x_0213_doublebyte_0xe7 = {
	0x40: [`\u8E47`].string() // U+8E47 <cjk>
	0x41: [`\u8E49`].string() // U+8E49 <cjk>
	0x42: [`\u8E4C`].string() // U+8E4C <cjk>
	0x43: [`\u8E50`].string() // U+8E50 <cjk>
	0x44: [`\u8E48`].string() // U+8E48 <cjk>
	0x45: [`\u8E59`].string() // U+8E59 <cjk>
	0x46: [`\u8E64`].string() // U+8E64 <cjk>
	0x47: [`\u8E60`].string() // U+8E60 <cjk>
	0x48: [`\u8E2A`].string() // U+8E2A <cjk>
	0x49: [`\u8E63`].string() // U+8E63 <cjk>
	0x4A: [`\u8E55`].string() // U+8E55 <cjk>
	0x4B: [`\u8E76`].string() // U+8E76 <cjk>
	0x4C: [`\u8E72`].string() // U+8E72 <cjk>
	0x4D: [`\u8E7C`].string() // U+8E7C <cjk>
	0x4E: [`\u8E81`].string() // U+8E81 <cjk>
	0x4F: [`\u8E87`].string() // U+8E87 <cjk>
	0x50: [`\u8E85`].string() // U+8E85 <cjk>
	0x51: [`\u8E84`].string() // U+8E84 <cjk>
	0x52: [`\u8E8B`].string() // U+8E8B <cjk>
	0x53: [`\u8E8A`].string() // U+8E8A <cjk>
	0x54: [`\u8E93`].string() // U+8E93 <cjk>
	0x55: [`\u8E91`].string() // U+8E91 <cjk>
	0x56: [`\u8E94`].string() // U+8E94 <cjk>
	0x57: [`\u8E99`].string() // U+8E99 <cjk>
	0x58: [`\u8EAA`].string() // U+8EAA <cjk>
	0x59: [`\u8EA1`].string() // U+8EA1 <cjk>
	0x5A: [`\u8EAC`].string() // U+8EAC <cjk>
	0x5B: [`\u8EB0`].string() // U+8EB0 <cjk>
	0x5C: [`\u8EC6`].string() // U+8EC6 <cjk>
	0x5D: [`\u8EB1`].string() // U+8EB1 <cjk>
	0x5E: [`\u8EBE`].string() // U+8EBE <cjk>
	0x5F: [`\u8EC5`].string() // U+8EC5 <cjk>
	0x60: [`\u8EC8`].string() // U+8EC8 <cjk>
	0x61: [`\u8ECB`].string() // U+8ECB <cjk>
	0x62: [`\u8EDB`].string() // U+8EDB <cjk>
	0x63: [`\u8EE3`].string() // U+8EE3 <cjk>
	0x64: [`\u8EFC`].string() // U+8EFC <cjk>
	0x65: [`\u8EFB`].string() // U+8EFB <cjk>
	0x66: [`\u8EEB`].string() // U+8EEB <cjk>
	0x67: [`\u8EFE`].string() // U+8EFE <cjk>
	0x68: [`\u8F0A`].string() // U+8F0A <cjk>
	0x69: [`\u8F05`].string() // U+8F05 <cjk>
	0x6A: [`\u8F15`].string() // U+8F15 <cjk>
	0x6B: [`\u8F12`].string() // U+8F12 <cjk>
	0x6C: [`\u8F19`].string() // U+8F19 <cjk>
	0x6D: [`\u8F13`].string() // U+8F13 <cjk>
	0x6E: [`\u8F1C`].string() // U+8F1C <cjk>
	0x6F: [`\u8F1F`].string() // U+8F1F <cjk>
	0x70: [`\u8F1B`].string() // U+8F1B <cjk>
	0x71: [`\u8F0C`].string() // U+8F0C <cjk>
	0x72: [`\u8F26`].string() // U+8F26 <cjk>
	0x73: [`\u8F33`].string() // U+8F33 <cjk>
	0x74: [`\u8F3B`].string() // U+8F3B <cjk>
	0x75: [`\u8F39`].string() // U+8F39 <cjk>
	0x76: [`\u8F45`].string() // U+8F45 <cjk>
	0x77: [`\u8F42`].string() // U+8F42 <cjk>
	0x78: [`\u8F3E`].string() // U+8F3E <cjk>
	0x79: [`\u8F4C`].string() // U+8F4C <cjk>
	0x7A: [`\u8F49`].string() // U+8F49 <cjk>
	0x7B: [`\u8F46`].string() // U+8F46 <cjk>
	0x7C: [`\u8F4E`].string() // U+8F4E <cjk>
	0x7D: [`\u8F57`].string() // U+8F57 <cjk>
	0x7E: [`\u8F5C`].string() // U+8F5C <cjk>
	0x80: [`\u8F62`].string() // U+8F62 <cjk>
	0x81: [`\u8F63`].string() // U+8F63 <cjk>
	0x82: [`\u8F64`].string() // U+8F64 <cjk>
	0x83: [`\u8F9C`].string() // U+8F9C <cjk>
	0x84: [`\u8F9F`].string() // U+8F9F <cjk>
	0x85: [`\u8FA3`].string() // U+8FA3 <cjk>
	0x86: [`\u8FAD`].string() // U+8FAD <cjk>
	0x87: [`\u8FAF`].string() // U+8FAF <cjk>
	0x88: [`\u8FB7`].string() // U+8FB7 <cjk>
	0x89: [`\u8FDA`].string() // U+8FDA <cjk>
	0x8A: [`\u8FE5`].string() // U+8FE5 <cjk>
	0x8B: [`\u8FE2`].string() // U+8FE2 <cjk>
	0x8C: [`\u8FEA`].string() // U+8FEA <cjk>
	0x8D: [`\u8FEF`].string() // U+8FEF <cjk>
	0x8E: [`\u9087`].string() // U+9087 <cjk>
	0x8F: [`\u8FF4`].string() // U+8FF4 <cjk>
	0x90: [`\u9005`].string() // U+9005 <cjk>
	0x91: [`\u8FF9`].string() // U+8FF9 <cjk>
	0x92: [`\u8FFA`].string() // U+8FFA <cjk>
	0x93: [`\u9011`].string() // U+9011 <cjk>
	0x94: [`\u9015`].string() // U+9015 <cjk>
	0x95: [`\u9021`].string() // U+9021 <cjk>
	0x96: [`\u900D`].string() // U+900D <cjk>
	0x97: [`\u901E`].string() // U+901E <cjk>
	0x98: [`\u9016`].string() // U+9016 <cjk>
	0x99: [`\u900B`].string() // U+900B <cjk>
	0x9A: [`\u9027`].string() // U+9027 <cjk>
	0x9B: [`\u9036`].string() // U+9036 <cjk>
	0x9C: [`\u9035`].string() // U+9035 <cjk>
	0x9D: [`\u9039`].string() // U+9039 <cjk>
	0x9E: [`\u8FF8`].string() // U+8FF8 <cjk>
	0x9F: [`\u904F`].string() // U+904F <cjk>
	0xA0: [`\u9050`].string() // U+9050 <cjk>
	0xA1: [`\u9051`].string() // U+9051 <cjk>
	0xA2: [`\u9052`].string() // U+9052 <cjk>
	0xA3: [`\u900E`].string() // U+900E <cjk>
	0xA4: [`\u9049`].string() // U+9049 <cjk>
	0xA5: [`\u903E`].string() // U+903E <cjk>
	0xA6: [`\u9056`].string() // U+9056 <cjk>
	0xA7: [`\u9058`].string() // U+9058 <cjk>
	0xA8: [`\u905E`].string() // U+905E <cjk>
	0xA9: [`\u9068`].string() // U+9068 <cjk>
	0xAA: [`\u906F`].string() // U+906F <cjk>
	0xAB: [`\u9076`].string() // U+9076 <cjk>
	0xAC: [`\u96A8`].string() // U+96A8 <cjk>
	0xAD: [`\u9072`].string() // U+9072 <cjk>
	0xAE: [`\u9082`].string() // U+9082 <cjk>
	0xAF: [`\u907D`].string() // U+907D <cjk>
	0xB0: [`\u9081`].string() // U+9081 <cjk>
	0xB1: [`\u9080`].string() // U+9080 <cjk>
	0xB2: [`\u908A`].string() // U+908A <cjk>
	0xB3: [`\u9089`].string() // U+9089 <cjk>
	0xB4: [`\u908F`].string() // U+908F <cjk>
	0xB5: [`\u90A8`].string() // U+90A8 <cjk>
	0xB6: [`\u90AF`].string() // U+90AF <cjk>
	0xB7: [`\u90B1`].string() // U+90B1 <cjk>
	0xB8: [`\u90B5`].string() // U+90B5 <cjk>
	0xB9: [`\u90E2`].string() // U+90E2 <cjk>
	0xBA: [`\u90E4`].string() // U+90E4 <cjk>
	0xBB: [`\u6248`].string() // U+6248 <cjk>
	0xBC: [`\u90DB`].string() // U+90DB <cjk>
	0xBD: [`\u9102`].string() // U+9102 <cjk>
	0xBE: [`\u9112`].string() // U+9112 <cjk>
	0xBF: [`\u9119`].string() // U+9119 <cjk>
	0xC0: [`\u9132`].string() // U+9132 <cjk>
	0xC1: [`\u9130`].string() // U+9130 <cjk>
	0xC2: [`\u914A`].string() // U+914A <cjk>
	0xC3: [`\u9156`].string() // U+9156 <cjk>
	0xC4: [`\u9158`].string() // U+9158 <cjk>
	0xC5: [`\u9163`].string() // U+9163 <cjk>
	0xC6: [`\u9165`].string() // U+9165 <cjk>
	0xC7: [`\u9169`].string() // U+9169 <cjk>
	0xC8: [`\u9173`].string() // U+9173 <cjk>
	0xC9: [`\u9172`].string() // U+9172 <cjk>
	0xCA: [`\u918B`].string() // U+918B <cjk>
	0xCB: [`\u9189`].string() // U+9189 <cjk>
	0xCC: [`\u9182`].string() // U+9182 <cjk>
	0xCD: [`\u91A2`].string() // U+91A2 <cjk>
	0xCE: [`\u91AB`].string() // U+91AB <cjk>
	0xCF: [`\u91AF`].string() // U+91AF <cjk>
	0xD0: [`\u91AA`].string() // U+91AA <cjk>
	0xD1: [`\u91B5`].string() // U+91B5 <cjk>
	0xD2: [`\u91B4`].string() // U+91B4 <cjk>
	0xD3: [`\u91BA`].string() // U+91BA <cjk>
	0xD4: [`\u91C0`].string() // U+91C0 <cjk>
	0xD5: [`\u91C1`].string() // U+91C1 <cjk>
	0xD6: [`\u91C9`].string() // U+91C9 <cjk>
	0xD7: [`\u91CB`].string() // U+91CB <cjk>
	0xD8: [`\u91D0`].string() // U+91D0 <cjk>
	0xD9: [`\u91D6`].string() // U+91D6 <cjk>
	0xDA: [`\u91DF`].string() // U+91DF <cjk>
	0xDB: [`\u91E1`].string() // U+91E1 <cjk>
	0xDC: [`\u91DB`].string() // U+91DB <cjk>
	0xDD: [`\u91FC`].string() // U+91FC <cjk>
	0xDE: [`\u91F5`].string() // U+91F5 <cjk>
	0xDF: [`\u91F6`].string() // U+91F6 <cjk>
	0xE0: [`\u921E`].string() // U+921E <cjk>
	0xE1: [`\u91FF`].string() // U+91FF <cjk>
	0xE2: [`\u9214`].string() // U+9214 <cjk>
	0xE3: [`\u922C`].string() // U+922C <cjk>
	0xE4: [`\u9215`].string() // U+9215 <cjk>
	0xE5: [`\u9211`].string() // U+9211 <cjk>
	0xE6: [`\u925E`].string() // U+925E <cjk>
	0xE7: [`\u9257`].string() // U+9257 <cjk>
	0xE8: [`\u9245`].string() // U+9245 <cjk>
	0xE9: [`\u9249`].string() // U+9249 <cjk>
	0xEA: [`\u9264`].string() // U+9264 <cjk>
	0xEB: [`\u9248`].string() // U+9248 <cjk>
	0xEC: [`\u9295`].string() // U+9295 <cjk>
	0xED: [`\u923F`].string() // U+923F <cjk>
	0xEE: [`\u924B`].string() // U+924B <cjk>
	0xEF: [`\u9250`].string() // U+9250 <cjk>
	0xF0: [`\u929C`].string() // U+929C <cjk>
	0xF1: [`\u9296`].string() // U+9296 <cjk>
	0xF2: [`\u9293`].string() // U+9293 <cjk>
	0xF3: [`\u929B`].string() // U+929B <cjk>
	0xF4: [`\u925A`].string() // U+925A <cjk>
	0xF5: [`\u92CF`].string() // U+92CF <cjk>
	0xF6: [`\u92B9`].string() // U+92B9 <cjk>
	0xF7: [`\u92B7`].string() // U+92B7 <cjk>
	0xF8: [`\u92E9`].string() // U+92E9 <cjk>
	0xF9: [`\u930F`].string() // U+930F <cjk>
	0xFA: [`\u92FA`].string() // U+92FA <cjk>
	0xFB: [`\u9344`].string() // U+9344 <cjk>
	0xFC: [`\u932E`].string() // U+932E <cjk>
}

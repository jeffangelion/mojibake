module mojibake

const jis_x_0213_doublebyte_0xee = {
	0x40: [`\u83D1`].string() // U+83D1 <cjk>
	0x41: [`\u83E1`].string() // U+83E1 <cjk>
	0x42: [`\u83EA`].string() // U+83EA <cjk>
	0x43: [`\u8401`].string() // U+8401 <cjk>
	0x44: [`\u8406`].string() // U+8406 <cjk>
	0x45: [`\u840A`].string() // U+840A <cjk>
	0x46: [`\uFA5F`].string() // U+FA5F CJK COMPATIBILITY IDEOGRAPH-FA5F
	0x47: [`\u8448`].string() // U+8448 <cjk>
	0x48: [`\u845F`].string() // U+845F <cjk>
	0x49: [`\u8470`].string() // U+8470 <cjk>
	0x4A: [`\u8473`].string() // U+8473 <cjk>
	0x4B: [`\u8485`].string() // U+8485 <cjk>
	0x4C: [`\u849E`].string() // U+849E <cjk>
	0x4D: [`\u84AF`].string() // U+84AF <cjk>
	0x4E: [`\u84B4`].string() // U+84B4 <cjk>
	0x4F: [`\u84BA`].string() // U+84BA <cjk>
	0x50: [`\u84C0`].string() // U+84C0 <cjk>
	0x51: [`\u84C2`].string() // U+84C2 <cjk>
	0x52: utf32_to_str(0x26E40) // U+26E40 <cjk>
	0x53: [`\u8532`].string() // U+8532 <cjk>
	0x54: [`\u851E`].string() // U+851E <cjk>
	0x55: [`\u8523`].string() // U+8523 <cjk>
	0x56: [`\u852F`].string() // U+852F <cjk>
	0x57: [`\u8559`].string() // U+8559 <cjk>
	0x58: [`\u8564`].string() // U+8564 <cjk>
	0x59: [`\uFA1F`].string() // U+FA1F CJK COMPATIBILITY IDEOGRAPH-FA1F
	0x5A: [`\u85AD`].string() // U+85AD <cjk>
	0x5B: [`\u857A`].string() // U+857A <cjk>
	0x5C: [`\u858C`].string() // U+858C <cjk>
	0x5D: [`\u858F`].string() // U+858F <cjk>
	0x5E: [`\u85A2`].string() // U+85A2 <cjk>
	0x5F: [`\u85B0`].string() // U+85B0 <cjk>
	0x60: [`\u85CB`].string() // U+85CB <cjk>
	0x61: [`\u85CE`].string() // U+85CE <cjk>
	0x62: [`\u85ED`].string() // U+85ED <cjk>
	0x63: [`\u8612`].string() // U+8612 <cjk>
	0x64: [`\u85FF`].string() // U+85FF <cjk>
	0x65: [`\u8604`].string() // U+8604 <cjk>
	0x66: [`\u8605`].string() // U+8605 <cjk>
	0x67: [`\u8610`].string() // U+8610 <cjk>
	0x68: utf32_to_str(0x270F4) // U+270F4 <cjk>
	0x69: [`\u8618`].string() // U+8618 <cjk>
	0x6A: [`\u8629`].string() // U+8629 <cjk>
	0x6B: [`\u8638`].string() // U+8638 <cjk>
	0x6C: [`\u8657`].string() // U+8657 <cjk>
	0x6D: [`\u865B`].string() // U+865B <cjk>
	0x6E: [`\uF936`].string() // U+F936 CJK COMPATIBILITY IDEOGRAPH-F936
	0x6F: [`\u8662`].string() // U+8662 <cjk>
	0x70: [`\u459D`].string() // U+459D <cjk>
	0x71: [`\u866C`].string() // U+866C <cjk>
	0x72: [`\u8675`].string() // U+8675 <cjk>
	0x73: [`\u8698`].string() // U+8698 <cjk>
	0x74: [`\u86B8`].string() // U+86B8 <cjk>
	0x75: [`\u86FA`].string() // U+86FA <cjk>
	0x76: [`\u86FC`].string() // U+86FC <cjk>
	0x77: [`\u86FD`].string() // U+86FD <cjk>
	0x78: [`\u870B`].string() // U+870B <cjk>
	0x79: [`\u8771`].string() // U+8771 <cjk>
	0x7A: [`\u8787`].string() // U+8787 <cjk>
	0x7B: [`\u8788`].string() // U+8788 <cjk>
	0x7C: [`\u87AC`].string() // U+87AC <cjk>
	0x7D: [`\u87AD`].string() // U+87AD <cjk>
	0x7E: [`\u87B5`].string() // U+87B5 <cjk>
	0x80: [`\u45EA`].string() // U+45EA <cjk>
	0x81: [`\u87D6`].string() // U+87D6 <cjk>
	0x82: [`\u87EC`].string() // U+87EC <cjk>
	0x83: [`\u8806`].string() // U+8806 <cjk>
	0x84: [`\u880A`].string() // U+880A <cjk>
	0x85: [`\u8810`].string() // U+8810 <cjk>
	0x86: [`\u8814`].string() // U+8814 <cjk>
	0x87: [`\u881F`].string() // U+881F <cjk>
	0x88: [`\u8898`].string() // U+8898 <cjk>
	0x89: [`\u88AA`].string() // U+88AA <cjk>
	0x8A: [`\u88CA`].string() // U+88CA <cjk>
	0x8B: [`\u88CE`].string() // U+88CE <cjk>
	0x8C: utf32_to_str(0x27684) // U+27684 <cjk>
	0x8D: [`\u88F5`].string() // U+88F5 <cjk>
	0x8E: [`\u891C`].string() // U+891C <cjk>
	0x8F: [`\uFA60`].string() // U+FA60 CJK COMPATIBILITY IDEOGRAPH-FA60
	0x90: [`\u8918`].string() // U+8918 <cjk>
	0x91: [`\u8919`].string() // U+8919 <cjk>
	0x92: [`\u891A`].string() // U+891A <cjk>
	0x93: [`\u8927`].string() // U+8927 <cjk>
	0x94: [`\u8930`].string() // U+8930 <cjk>
	0x95: [`\u8932`].string() // U+8932 <cjk>
	0x96: [`\u8939`].string() // U+8939 <cjk>
	0x97: [`\u8940`].string() // U+8940 <cjk>
	0x98: [`\u8994`].string() // U+8994 <cjk>
	0x99: [`\uFA61`].string() // U+FA61 CJK COMPATIBILITY IDEOGRAPH-FA61
	0x9A: [`\u89D4`].string() // U+89D4 <cjk>
	0x9B: [`\u89E5`].string() // U+89E5 <cjk>
	0x9C: [`\u89F6`].string() // U+89F6 <cjk>
	0x9D: [`\u8A12`].string() // U+8A12 <cjk>
	0x9E: [`\u8A15`].string() // U+8A15 <cjk>
	0x9F: [`\u8A22`].string() // U+8A22 <cjk>
	0xA0: [`\u8A37`].string() // U+8A37 <cjk>
	0xA1: [`\u8A47`].string() // U+8A47 <cjk>
	0xA2: [`\u8A4E`].string() // U+8A4E <cjk>
	0xA3: [`\u8A5D`].string() // U+8A5D <cjk>
	0xA4: [`\u8A61`].string() // U+8A61 <cjk>
	0xA5: [`\u8A75`].string() // U+8A75 <cjk>
	0xA6: [`\u8A79`].string() // U+8A79 <cjk>
	0xA7: [`\u8AA7`].string() // U+8AA7 <cjk>
	0xA8: [`\u8AD0`].string() // U+8AD0 <cjk>
	0xA9: [`\u8ADF`].string() // U+8ADF <cjk>
	0xAA: [`\u8AF4`].string() // U+8AF4 <cjk>
	0xAB: [`\u8AF6`].string() // U+8AF6 <cjk>
	0xAC: [`\uFA22`].string() // U+FA22 CJK COMPATIBILITY IDEOGRAPH-FA22
	0xAD: [`\uFA62`].string() // U+FA62 CJK COMPATIBILITY IDEOGRAPH-FA62
	0xAE: [`\uFA63`].string() // U+FA63 CJK COMPATIBILITY IDEOGRAPH-FA63
	0xAF: [`\u8B46`].string() // U+8B46 <cjk>
	0xB0: [`\u8B54`].string() // U+8B54 <cjk>
	0xB1: [`\u8B59`].string() // U+8B59 <cjk>
	0xB2: [`\u8B69`].string() // U+8B69 <cjk>
	0xB3: [`\u8B9D`].string() // U+8B9D <cjk>
	0xB4: [`\u8C49`].string() // U+8C49 <cjk>
	0xB5: [`\u8C68`].string() // U+8C68 <cjk>
	0xB6: [`\uFA64`].string() // U+FA64 CJK COMPATIBILITY IDEOGRAPH-FA64
	0xB7: [`\u8CE1`].string() // U+8CE1 <cjk>
	0xB8: [`\u8CF4`].string() // U+8CF4 <cjk>
	0xB9: [`\u8CF8`].string() // U+8CF8 <cjk>
	0xBA: [`\u8CFE`].string() // U+8CFE <cjk>
	0xBB: [`\uFA65`].string() // U+FA65 CJK COMPATIBILITY IDEOGRAPH-FA65
	0xBC: [`\u8D12`].string() // U+8D12 <cjk>
	0xBD: [`\u8D1B`].string() // U+8D1B <cjk>
	0xBE: [`\u8DAF`].string() // U+8DAF <cjk>
	0xBF: [`\u8DCE`].string() // U+8DCE <cjk>
	0xC0: [`\u8DD1`].string() // U+8DD1 <cjk>
	0xC1: [`\u8DD7`].string() // U+8DD7 <cjk>
	0xC2: [`\u8E20`].string() // U+8E20 <cjk>
	0xC3: [`\u8E23`].string() // U+8E23 <cjk>
	0xC4: [`\u8E3D`].string() // U+8E3D <cjk>
	0xC5: [`\u8E70`].string() // U+8E70 <cjk>
	0xC6: [`\u8E7B`].string() // U+8E7B <cjk>
	0xC7: utf32_to_str(0x28277) // U+28277 <cjk>
	0xC8: [`\u8EC0`].string() // U+8EC0 <cjk>
	0xC9: [`\u4844`].string() // U+4844 <cjk>
	0xCA: [`\u8EFA`].string() // U+8EFA <cjk>
	0xCB: [`\u8F1E`].string() // U+8F1E <cjk>
	0xCC: [`\u8F2D`].string() // U+8F2D <cjk>
	0xCD: [`\u8F36`].string() // U+8F36 <cjk>
	0xCE: [`\u8F54`].string() // U+8F54 <cjk>
	0xCF: utf32_to_str(0x283CD) // U+283CD <cjk>
	0xD0: [`\u8FA6`].string() // U+8FA6 <cjk>
	0xD1: [`\u8FB5`].string() // U+8FB5 <cjk>
	0xD2: [`\u8FE4`].string() // U+8FE4 <cjk>
	0xD3: [`\u8FE8`].string() // U+8FE8 <cjk>
	0xD4: [`\u8FEE`].string() // U+8FEE <cjk>
	0xD5: [`\u9008`].string() // U+9008 <cjk>
	0xD6: [`\u902D`].string() // U+902D <cjk>
	0xD7: [`\uFA67`].string() // U+FA67 CJK COMPATIBILITY IDEOGRAPH-FA67
	0xD8: [`\u9088`].string() // U+9088 <cjk>
	0xD9: [`\u9095`].string() // U+9095 <cjk>
	0xDA: [`\u9097`].string() // U+9097 <cjk>
	0xDB: [`\u9099`].string() // U+9099 <cjk>
	0xDC: [`\u909B`].string() // U+909B <cjk>
	0xDD: [`\u90A2`].string() // U+90A2 <cjk>
	0xDE: [`\u90B3`].string() // U+90B3 <cjk>
	0xDF: [`\u90BE`].string() // U+90BE <cjk>
	0xE0: [`\u90C4`].string() // U+90C4 <cjk>
	0xE1: [`\u90C5`].string() // U+90C5 <cjk>
	0xE2: [`\u90C7`].string() // U+90C7 <cjk>
	0xE3: [`\u90D7`].string() // U+90D7 <cjk>
	0xE4: [`\u90DD`].string() // U+90DD <cjk>
	0xE5: [`\u90DE`].string() // U+90DE <cjk>
	0xE6: [`\u90EF`].string() // U+90EF <cjk>
	0xE7: [`\u90F4`].string() // U+90F4 <cjk>
	0xE8: [`\uFA26`].string() // U+FA26 CJK COMPATIBILITY IDEOGRAPH-FA26
	0xE9: [`\u9114`].string() // U+9114 <cjk>
	0xEA: [`\u9115`].string() // U+9115 <cjk>
	0xEB: [`\u9116`].string() // U+9116 <cjk>
	0xEC: [`\u9122`].string() // U+9122 <cjk>
	0xED: [`\u9123`].string() // U+9123 <cjk>
	0xEE: [`\u9127`].string() // U+9127 <cjk>
	0xEF: [`\u912F`].string() // U+912F <cjk>
	0xF0: [`\u9131`].string() // U+9131 <cjk>
	0xF1: [`\u9134`].string() // U+9134 <cjk>
	0xF2: [`\u913D`].string() // U+913D <cjk>
	0xF3: [`\u9148`].string() // U+9148 <cjk>
	0xF4: [`\u915B`].string() // U+915B <cjk>
	0xF5: [`\u9183`].string() // U+9183 <cjk>
	0xF6: [`\u919E`].string() // U+919E <cjk>
	0xF7: [`\u91AC`].string() // U+91AC <cjk>
	0xF8: [`\u91B1`].string() // U+91B1 <cjk>
	0xF9: [`\u91BC`].string() // U+91BC <cjk>
	0xFA: [`\u91D7`].string() // U+91D7 <cjk>
	0xFB: [`\u91FB`].string() // U+91FB <cjk>
	0xFC: [`\u91E4`].string() // U+91E4 <cjk>
}

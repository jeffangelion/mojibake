module mojibake

const jis_x_0213_doublebyte_0x81 = {
	0x40: [`\u3000`].string() // U+3000 IDEOGRAPHIC SPACE
	0x41: [`\u3001`].string() // U+3001 IDEOGRAPHIC COMMA
	0x42: [`\u3002`].string() // U+3002 IDEOGRAPHIC FULL STOP
	0x43: [`\uFF0C`].string() // U+FF0C FULLWIDTH COMMA
	0x44: [`\uFF0E`].string() // U+FF0E FULLWIDTH FULL STOP
	0x45: [`\u30FB`].string() // U+30FB KATAKANA MIDDLE DOT
	0x46: [`\uFF1A`].string() // U+FF1A FULLWIDTH COLON
	0x47: [`\uFF1B`].string() // U+FF1B FULLWIDTH SEMICOLON
	0x48: [`\uFF1F`].string() // U+FF1F FULLWIDTH QUESTION MARK
	0x49: [`\uFF01`].string() // U+FF01 FULLWIDTH EXCLAMATION MARK
	0x4A: [`\u309B`].string() // U+309B KATAKANA-HIRAGANA VOICED SOUND MARK
	0x4B: [`\u309C`].string() // U+309C KATAKANA-HIRAGANA SEMI-VOICED SOUND MARK
	0x4C: [`\u00B4`].string() // U+00B4 ACUTE ACCENT
	0x4D: [`\uFF40`].string() // U+FF40 FULLWIDTH GRAVE ACCENT
	0x4E: [`\u00A8`].string() // U+00A8 DIAERESIS
	0x4F: [`\uFF3E`].string() // U+FF3E FULLWIDTH CIRCUMFLEX ACCENT
	0x50: [`\uFFE3`].string() // U+FFE3 FULLWIDTH MACRON 
	0x51: [`\uFF3F`].string() // U+FF3F FULLWIDTH LOW LINE
	0x52: [`\u30FD`].string() // U+30FD KATAKANA ITERATION MARK
	0x53: [`\u30FE`].string() // U+30FE KATAKANA VOICED ITERATION MARK
	0x54: [`\u309D`].string() // U+309D HIRAGANA ITERATION MARK
	0x55: [`\u309E`].string() // U+309E HIRAGANA VOICED ITERATION MARK
	0x56: [`\u3003`].string() // U+3003 DITTO MARK
	0x57: [`\u4EDD`].string() // U+4EDD <cjk>
	0x58: [`\u3005`].string() // U+3005 IDEOGRAPHIC ITERATION MARK
	0x59: [`\u3006`].string() // U+3006 IDEOGRAPHIC CLOSING MARK
	0x5A: [`\u3007`].string() // U+3007 IDEOGRAPHIC NUMBER ZERO
	0x5B: [`\u30FC`].string() // U+30FC KATAKANA-HIRAGANA PROLONGED SOUND MARK
	0x5C: [`\u2014`].string() // U+2014 EM DASH
	0x5D: [`\u2010`].string() // U+2010 HYPHEN
	0x5E: [`\uFF0F`].string() // U+FF0F FULLWIDTH SOLIDUS
	0x5F: [`\u005C`].string() // U+005C REVERSE SOLIDUS
	0x60: [`\u301C`].string() // U+301C WAVE DASH
	0x61: [`\u2016`].string() // U+2016 DOUBLE VERTICAL LINE
	0x62: [`\uFF5C`].string() // U+FF5C FULLWIDTH VERTICAL LINE
	0x63: [`\u2026`].string() // U+2026 HORIZONTAL ELLIPSIS
	0x64: [`\u2025`].string() // U+2025 TWO DOT LEADER
	0x65: [`\u2018`].string() // U+2018 LEFT SINGLE QUOTATION MARK
	0x66: [`\u2019`].string() // U+2019 RIGHT SINGLE QUOTATION MARK
	0x67: [`\u201C`].string() // U+201C LEFT DOUBLE QUOTATION MARK
	0x68: [`\u201D`].string() // U+201D RIGHT DOUBLE QUOTATION MARK
	0x69: [`\uFF08`].string() // U+FF08 FULLWIDTH LEFT PARENTHESIS
	0x6A: [`\uFF09`].string() // U+FF09 FULLWIDTH RIGHT PARENTHESIS
	0x6B: [`\u3014`].string() // U+3014 LEFT TORTOISE SHELL BRACKET
	0x6C: [`\u3015`].string() // U+3015 RIGHT TORTOISE SHELL BRACKET
	0x6D: [`\uFF3B`].string() // U+FF3B FULLWIDTH LEFT SQUARE BRACKET
	0x6E: [`\uFF3D`].string() // U+FF3D FULLWIDTH RIGHT SQUARE BRACKET
	0x6F: [`\uFF5B`].string() // U+FF5B FULLWIDTH LEFT CURLY BRACKET
	0x70: [`\uFF5D`].string() // U+FF5D FULLWIDTH RIGHT CURLY BRACKET
	0x71: [`\u3008`].string() // U+3008 LEFT ANGLE BRACKET
	0x72: [`\u3009`].string() // U+3009 RIGHT ANGLE BRACKET
	0x73: [`\u300A`].string() // U+300A LEFT DOUBLE ANGLE BRACKET
	0x74: [`\u300B`].string() // U+300B RIGHT DOUBLE ANGLE BRACKET
	0x75: [`\u300C`].string() // U+300C LEFT CORNER BRACKET
	0x76: [`\u300D`].string() // U+300D RIGHT CORNER BRACKET
	0x77: [`\u300E`].string() // U+300E LEFT WHITE CORNER BRACKET
	0x78: [`\u300F`].string() // U+300F RIGHT WHITE CORNER BRACKET
	0x79: [`\u3010`].string() // U+3010 LEFT BLACK LENTICULAR BRACKET
	0x7A: [`\u3011`].string() // U+3011 RIGHT BLACK LENTICULAR BRACKET
	0x7B: [`\uFF0B`].string() // U+FF0B FULLWIDTH PLUS SIGN
	0x7C: [`\u2212`].string() // U+2212 MINUS SIGN
	0x7D: [`\u00B1`].string() // U+00B1 PLUS-MINUS SIGN
	0x7E: [`\u00D7`].string() // U+00D7 MULTIPLICATION SIGN
	0x80: [`\u00F7`].string() // U+00F7 DIVISION SIGN
	0x81: [`\uFF1D`].string() // U+FF1D FULLWIDTH EQUALS SIGN
	0x82: [`\u2260`].string() // U+2260 NOT EQUAL TO
	0x83: [`\uFF1C`].string() // U+FF1C FULLWIDTH LESS-THAN SIGN
	0x84: [`\uFF1E`].string() // U+FF1E FULLWIDTH GREATER-THAN SIGN
	0x85: [`\u2266`].string() // U+2266 LESS-THAN OVER EQUAL TO
	0x86: [`\u2267`].string() // U+2267 GREATER-THAN OVER EQUAL TO
	0x87: [`\u221E`].string() // U+221E INFINITY
	0x88: [`\u2234`].string() // U+2234 THEREFORE
	0x89: [`\u2642`].string() // U+2642 MALE SIGN
	0x8A: [`\u2640`].string() // U+2640 FEMALE SIGN
	0x8B: [`\u00B0`].string() // U+00B0 DEGREE SIGN
	0x8C: [`\u2032`].string() // U+2032 PRIME
	0x8D: [`\u2033`].string() // U+2033 DOUBLE PRIME
	0x8E: [`\u2103`].string() // U+2103 DEGREE CELSIUS
	0x8F: [`\uFFE5`].string() // U+FFE5 FULLWIDTH YEN SIGN
	0x90: [`\uFF04`].string() // U+FF04 FULLWIDTH DOLLAR SIGN
	0x91: [`\u00A2`].string() // U+00A2 CENT SIGN
	0x92: [`\u00A3`].string() // U+00A3 POUND SIGN
	0x93: [`\uFF05`].string() // U+FF05 FULLWIDTH PERCENT SIGN
	0x94: [`\uFF03`].string() // U+FF03 FULLWIDTH NUMBER SIGN
	0x95: [`\uFF06`].string() // U+FF06 FULLWIDTH AMPERSAND
	0x96: [`\uFF0A`].string() // U+FF0A FULLWIDTH ASTERISK
	0x97: [`\uFF20`].string() // U+FF20 FULLWIDTH COMMERCIAL AT
	0x98: [`\u00A7`].string() // U+00A7 SECTION SIGN
	0x99: [`\u2606`].string() // U+2606 WHITE STAR
	0x9A: [`\u2605`].string() // U+2605 BLACK STAR
	0x9B: [`\u25CB`].string() // U+25CB WHITE CIRCLE
	0x9C: [`\u25CF`].string() // U+25CF BLACK CIRCLE
	0x9D: [`\u25CE`].string() // U+25CE BULLSEYE
	0x9E: [`\u25C7`].string() // U+25C7 WHITE DIAMOND
	0x9F: [`\u25C6`].string() // U+25C6 BLACK DIAMOND
	0xA0: [`\u25A1`].string() // U+25A1 WHITE SQUARE
	0xA1: [`\u25A0`].string() // U+25A0 BLACK SQUARE
	0xA2: [`\u25B3`].string() // U+25B3 WHITE UP-POINTING TRIANGLE
	0xA3: [`\u25B2`].string() // U+25B2 BLACK UP-POINTING TRIANGLE
	0xA4: [`\u25BD`].string() // U+25BD WHITE DOWN-POINTING TRIANGLE
	0xA5: [`\u25BC`].string() // U+25BC BLACK DOWN-POINTING TRIANGLE
	0xA6: [`\u203B`].string() // U+203B REFERENCE MARK
	0xA7: [`\u3012`].string() // U+3012 POSTAL MARK
	0xA8: [`\u2192`].string() // U+2192 RIGHTWARDS ARROW
	0xA9: [`\u2190`].string() // U+2190 LEFTWARDS ARROW
	0xAA: [`\u2191`].string() // U+2191 UPWARDS ARROW
	0xAB: [`\u2193`].string() // U+2193 DOWNWARDS ARROW
	0xAC: [`\u3013`].string() // U+3013 GETA MARK
	0xAD: [`\uFF07`].string() // U+FF07 FULLWIDTH APOSTROPHE
	0xAE: [`\uFF02`].string() // U+FF02 FULLWIDTH QUOTATION MARK
	0xAF: [`\uFF0D`].string() // U+FF0D FULLWIDTH HYPHEN-MINUS
	0xB0: [`\u007E`].string() // U+007E TILDE
	0xB1: [`\u3033`].string() // U+3033 VERTICAL KANA REPEAT MARK UPPER HALF
	0xB2: [`\u3034`].string() // U+3034 VERTICAL KANA REPEAT WITH VOICED SOUND MARK UPPER HALF
	0xB3: [`\u3035`].string() // U+3035 VERTICAL KANA REPEAT MARK LOWER HALF
	0xB4: [`\u303B`].string() // U+303B VERTICAL IDEOGRAPHIC ITERATION MARK
	0xB5: [`\u303C`].string() // U+303C MASU MARK
	0xB6: [`\u30FF`].string() // U+30FF KATAKANA DIGRAPH KOTO
	0xB7: [`\u309F`].string() // U+309F HIRAGANA DIGRAPH YORI
	0xB8: [`\u2208`].string() // U+2208 ELEMENT OF
	0xB9: [`\u220B`].string() // U+220B CONTAINS AS MEMBER
	0xBA: [`\u2286`].string() // U+2286 SUBSET OF OR EQUAL TO
	0xBB: [`\u2287`].string() // U+2287 SUPERSET OF OR EQUAL TO
	0xBC: [`\u2282`].string() // U+2282 SUBSET OF
	0xBD: [`\u2283`].string() // U+2283 SUPERSET OF
	0xBE: [`\u222A`].string() // U+222A UNION
	0xBF: [`\u2229`].string() // U+2229 INTERSECTION
	0xC0: [`\u2284`].string() // U+2284 NOT A SUBSET OF
	0xC1: [`\u2285`].string() // U+2285 NOT A SUPERSET OF
	0xC2: [`\u228A`].string() // U+228A SUBSET OF WITH NOT EQUAL TO
	0xC3: [`\u228B`].string() // U+228B SUPERSET OF WITH NOT EQUAL TO
	0xC4: [`\u2209`].string() // U+2209 NOT AN ELEMENT OF
	0xC5: [`\u2205`].string() // U+2205 EMPTY SET
	0xC6: [`\u2305`].string() // U+2305 PROJECTIVE
	0xC7: [`\u2306`].string() // U+2306 PERSPECTIVE
	0xC8: [`\u2227`].string() // U+2227 LOGICAL AND
	0xC9: [`\u2228`].string() // U+2228 LOGICAL OR
	0xCA: [`\u00AC`].string() // U+00AC NOT SIGN
	0xCB: [`\u21D2`].string() // U+21D2 RIGHTWARDS DOUBLE ARROW
	0xCC: [`\u21D4`].string() // U+21D4 LEFT RIGHT DOUBLE ARROW
	0xCD: [`\u2200`].string() // U+2200 FOR ALL
	0xCE: [`\u2203`].string() // U+2203 THERE EXISTS
	0xCF: [`\u2295`].string() // U+2295 CIRCLED PLUS
	0xD0: [`\u2296`].string() // U+2296 CIRCLED MINUS
	0xD1: [`\u2297`].string() // U+2297 CIRCLED TIMES
	0xD2: [`\u2225`].string() // U+2225 PARALLEL TO
	0xD3: [`\u2226`].string() // U+2226 NOT PARALLEL TO
	0xD4: [`\uFF5F`].string() // U+FF5F FULLWIDTH LEFT WHITE PARENTHESIS
	0xD5: [`\uFF60`].string() // U+FF60 FULLWIDTH RIGHT WHITE PARENTHESIS
	0xD6: [`\u3018`].string() // U+3018 LEFT WHITE TORTOISE SHELL BRACKET
	0xD7: [`\u3019`].string() // U+3019 RIGHT WHITE TORTOISE SHELL BRACKET
	0xD8: [`\u3016`].string() // U+3016 LEFT WHITE LENTICULAR BRACKET
	0xD9: [`\u3017`].string() // U+3017 RIGHT WHITE LENTICULAR BRACKET
	0xDA: [`\u2220`].string() // U+2220 ANGLE
	0xDB: [`\u22A5`].string() // U+22A5 UP TACK
	0xDC: [`\u2312`].string() // U+2312 ARC
	0xDD: [`\u2202`].string() // U+2202 PARTIAL DIFFERENTIAL
	0xDE: [`\u2207`].string() // U+2207 NABLA
	0xDF: [`\u2261`].string() // U+2261 IDENTICAL TO
	0xE0: [`\u2252`].string() // U+2252 APPROXIMATELY EQUAL TO OR THE IMAGE OF
	0xE1: [`\u226A`].string() // U+226A MUCH LESS-THAN
	0xE2: [`\u226B`].string() // U+226B MUCH GREATER-THAN
	0xE3: [`\u221A`].string() // U+221A SQUARE ROOT
	0xE4: [`\u223D`].string() // U+223D REVERSED TILDE 
	0xE5: [`\u221D`].string() // U+221D PROPORTIONAL TO
	0xE6: [`\u2235`].string() // U+2235 BECAUSE
	0xE7: [`\u222B`].string() // U+222B INTEGRAL
	0xE8: [`\u222C`].string() // U+222C DOUBLE INTEGRAL
	0xE9: [`\u2262`].string() // U+2262 NOT IDENTICAL TO
	0xEA: [`\u2243`].string() // U+2243 ASYMPTOTICALLY EQUAL TO
	0xEB: [`\u2245`].string() // U+2245 APPROXIMATELY EQUAL TO
	0xEC: [`\u2248`].string() // U+2248 ALMOST EQUAL TO
	0xED: [`\u2276`].string() // U+2276 LESS-THAN OR GREATER-THAN
	0xEE: [`\u2277`].string() // U+2277 GREATER-THAN OR LESS-THAN
	0xEF: [`\u2194`].string() // U+2194 LEFT RIGHT ARROW
	0xF0: [`\u212B`].string() // U+212B ANGSTROM SIGN
	0xF1: [`\u2030`].string() // U+2030 PER MILLE SIGN
	0xF2: [`\u266F`].string() // U+266F MUSIC SHARP SIGN
	0xF3: [`\u266D`].string() // U+266D MUSIC FLAT SIGN
	0xF4: [`\u266A`].string() // U+266A EIGHTH NOTE
	0xF5: [`\u2020`].string() // U+2020 DAGGER
	0xF6: [`\u2021`].string() // U+2021 DOUBLE DAGGER
	0xF7: [`\u00B6`].string() // U+00B6 PILCROW SIGN
	0xF8: [`\u266E`].string() // U+266E MUSIC NATURAL SIGN
	0xF9: [`\u266B`].string() // U+266B BEAMED EIGHTH NOTES
	0xFA: [`\u266C`].string() // U+266C BEAMED SIXTEENTH NOTES
	0xFB: [`\u2669`].string() // U+2669 QUARTER NOTE
	0xFC: [`\u25EF`].string() // U+25EF LARGE CIRCLE
}

module mojibake

const jis_x_0213_doublebyte_0xe4 = {
	0x40: [`\u968B`].string() // U+968B <cjk>
	0x41: [`\u8146`].string() // U+8146 <cjk>
	0x42: [`\u813E`].string() // U+813E <cjk>
	0x43: [`\u8153`].string() // U+8153 <cjk>
	0x44: [`\u8151`].string() // U+8151 <cjk>
	0x45: [`\u80FC`].string() // U+80FC <cjk>
	0x46: [`\u8171`].string() // U+8171 <cjk>
	0x47: [`\u816E`].string() // U+816E <cjk>
	0x48: [`\u8165`].string() // U+8165 <cjk>
	0x49: [`\u8166`].string() // U+8166 <cjk>
	0x4A: [`\u8174`].string() // U+8174 <cjk>
	0x4B: [`\u8183`].string() // U+8183 <cjk>
	0x4C: [`\u8188`].string() // U+8188 <cjk>
	0x4D: [`\u818A`].string() // U+818A <cjk>
	0x4E: [`\u8180`].string() // U+8180 <cjk>
	0x4F: [`\u8182`].string() // U+8182 <cjk>
	0x50: [`\u81A0`].string() // U+81A0 <cjk>
	0x51: [`\u8195`].string() // U+8195 <cjk>
	0x52: [`\u81A4`].string() // U+81A4 <cjk>
	0x53: [`\u81A3`].string() // U+81A3 <cjk>
	0x54: [`\u815F`].string() // U+815F <cjk>
	0x55: [`\u8193`].string() // U+8193 <cjk>
	0x56: [`\u81A9`].string() // U+81A9 <cjk>
	0x57: [`\u81B0`].string() // U+81B0 <cjk>
	0x58: [`\u81B5`].string() // U+81B5 <cjk>
	0x59: [`\u81BE`].string() // U+81BE <cjk>
	0x5A: [`\u81B8`].string() // U+81B8 <cjk>
	0x5B: [`\u81BD`].string() // U+81BD <cjk>
	0x5C: [`\u81C0`].string() // U+81C0 <cjk>
	0x5D: [`\u81C2`].string() // U+81C2 <cjk>
	0x5E: [`\u81BA`].string() // U+81BA <cjk>
	0x5F: [`\u81C9`].string() // U+81C9 <cjk>
	0x60: [`\u81CD`].string() // U+81CD <cjk>
	0x61: [`\u81D1`].string() // U+81D1 <cjk>
	0x62: [`\u81D9`].string() // U+81D9 <cjk>
	0x63: [`\u81D8`].string() // U+81D8 <cjk>
	0x64: [`\u81C8`].string() // U+81C8 <cjk>
	0x65: [`\u81DA`].string() // U+81DA <cjk>
	0x66: [`\u81DF`].string() // U+81DF <cjk>
	0x67: [`\u81E0`].string() // U+81E0 <cjk>
	0x68: [`\u81E7`].string() // U+81E7 <cjk>
	0x69: [`\u81FA`].string() // U+81FA <cjk>
	0x6A: [`\u81FB`].string() // U+81FB <cjk>
	0x6B: [`\u81FE`].string() // U+81FE <cjk>
	0x6C: [`\u8201`].string() // U+8201 <cjk>
	0x6D: [`\u8202`].string() // U+8202 <cjk>
	0x6E: [`\u8205`].string() // U+8205 <cjk>
	0x6F: [`\u8207`].string() // U+8207 <cjk>
	0x70: [`\u820A`].string() // U+820A <cjk>
	0x71: [`\u820D`].string() // U+820D <cjk>
	0x72: [`\u8210`].string() // U+8210 <cjk>
	0x73: [`\u8216`].string() // U+8216 <cjk>
	0x74: [`\u8229`].string() // U+8229 <cjk>
	0x75: [`\u822B`].string() // U+822B <cjk>
	0x76: [`\u8238`].string() // U+8238 <cjk>
	0x77: [`\u8233`].string() // U+8233 <cjk>
	0x78: [`\u8240`].string() // U+8240 <cjk>
	0x79: [`\u8259`].string() // U+8259 <cjk>
	0x7A: [`\u8258`].string() // U+8258 <cjk>
	0x7B: [`\u825D`].string() // U+825D <cjk>
	0x7C: [`\u825A`].string() // U+825A <cjk>
	0x7D: [`\u825F`].string() // U+825F <cjk>
	0x7E: [`\u8264`].string() // U+8264 <cjk>
	0x80: [`\u8262`].string() // U+8262 <cjk>
	0x81: [`\u8268`].string() // U+8268 <cjk>
	0x82: [`\u826A`].string() // U+826A <cjk>
	0x83: [`\u826B`].string() // U+826B <cjk>
	0x84: [`\u822E`].string() // U+822E <cjk>
	0x85: [`\u8271`].string() // U+8271 <cjk>
	0x86: [`\u8277`].string() // U+8277 <cjk>
	0x87: [`\u8278`].string() // U+8278 <cjk>
	0x88: [`\u827E`].string() // U+827E <cjk>
	0x89: [`\u828D`].string() // U+828D <cjk>
	0x8A: [`\u8292`].string() // U+8292 <cjk>
	0x8B: [`\u82AB`].string() // U+82AB <cjk>
	0x8C: [`\u829F`].string() // U+829F <cjk>
	0x8D: [`\u82BB`].string() // U+82BB <cjk>
	0x8E: [`\u82AC`].string() // U+82AC <cjk>
	0x8F: [`\u82E1`].string() // U+82E1 <cjk>
	0x90: [`\u82E3`].string() // U+82E3 <cjk>
	0x91: [`\u82DF`].string() // U+82DF <cjk>
	0x92: [`\u82D2`].string() // U+82D2 <cjk>
	0x93: [`\u82F4`].string() // U+82F4 <cjk>
	0x94: [`\u82F3`].string() // U+82F3 <cjk>
	0x95: [`\u82FA`].string() // U+82FA <cjk>
	0x96: [`\u8393`].string() // U+8393 <cjk>
	0x97: [`\u8303`].string() // U+8303 <cjk>
	0x98: [`\u82FB`].string() // U+82FB <cjk>
	0x99: [`\u82F9`].string() // U+82F9 <cjk>
	0x9A: [`\u82DE`].string() // U+82DE <cjk>
	0x9B: [`\u8306`].string() // U+8306 <cjk>
	0x9C: [`\u82DC`].string() // U+82DC <cjk>
	0x9D: [`\u8309`].string() // U+8309 <cjk>
	0x9E: [`\u82D9`].string() // U+82D9 <cjk>
	0x9F: [`\u8335`].string() // U+8335 <cjk>
	0xA0: [`\u8334`].string() // U+8334 <cjk>
	0xA1: [`\u8316`].string() // U+8316 <cjk>
	0xA2: [`\u8332`].string() // U+8332 <cjk>
	0xA3: [`\u8331`].string() // U+8331 <cjk>
	0xA4: [`\u8340`].string() // U+8340 <cjk>
	0xA5: [`\u8339`].string() // U+8339 <cjk>
	0xA6: [`\u8350`].string() // U+8350 <cjk>
	0xA7: [`\u8345`].string() // U+8345 <cjk>
	0xA8: [`\u832F`].string() // U+832F <cjk>
	0xA9: [`\u832B`].string() // U+832B <cjk>
	0xAA: [`\u8317`].string() // U+8317 <cjk>
	0xAB: [`\u8318`].string() // U+8318 <cjk>
	0xAC: [`\u8385`].string() // U+8385 <cjk>
	0xAD: [`\u839A`].string() // U+839A <cjk>
	0xAE: [`\u83AA`].string() // U+83AA <cjk>
	0xAF: [`\u839F`].string() // U+839F <cjk>
	0xB0: [`\u83A2`].string() // U+83A2 <cjk>
	0xB1: [`\u8396`].string() // U+8396 <cjk>
	0xB2: [`\u8323`].string() // U+8323 <cjk>
	0xB3: [`\u838E`].string() // U+838E <cjk>
	0xB4: [`\u8387`].string() // U+8387 <cjk>
	0xB5: [`\u838A`].string() // U+838A <cjk>
	0xB6: [`\u837C`].string() // U+837C <cjk>
	0xB7: [`\u83B5`].string() // U+83B5 <cjk>
	0xB8: [`\u8373`].string() // U+8373 <cjk>
	0xB9: [`\u8375`].string() // U+8375 <cjk>
	0xBA: [`\u83A0`].string() // U+83A0 <cjk>
	0xBB: [`\u8389`].string() // U+8389 <cjk>
	0xBC: [`\u83A8`].string() // U+83A8 <cjk>
	0xBD: [`\u83F4`].string() // U+83F4 <cjk>
	0xBE: [`\u8413`].string() // U+8413 <cjk>
	0xBF: [`\u83EB`].string() // U+83EB <cjk>
	0xC0: [`\u83CE`].string() // U+83CE <cjk>
	0xC1: [`\u83FD`].string() // U+83FD <cjk>
	0xC2: [`\u8403`].string() // U+8403 <cjk>
	0xC3: [`\u83D8`].string() // U+83D8 <cjk>
	0xC4: [`\u840B`].string() // U+840B <cjk>
	0xC5: [`\u83C1`].string() // U+83C1 <cjk>
	0xC6: [`\u83F7`].string() // U+83F7 <cjk>
	0xC7: [`\u8407`].string() // U+8407 <cjk>
	0xC8: [`\u83E0`].string() // U+83E0 <cjk>
	0xC9: [`\u83F2`].string() // U+83F2 <cjk>
	0xCA: [`\u840D`].string() // U+840D <cjk>
	0xCB: [`\u8422`].string() // U+8422 <cjk>
	0xCC: [`\u8420`].string() // U+8420 <cjk>
	0xCD: [`\u83BD`].string() // U+83BD <cjk>
	0xCE: [`\u8438`].string() // U+8438 <cjk>
	0xCF: [`\u8506`].string() // U+8506 <cjk>
	0xD0: [`\u83FB`].string() // U+83FB <cjk>
	0xD1: [`\u846D`].string() // U+846D <cjk>
	0xD2: [`\u842A`].string() // U+842A <cjk>
	0xD3: [`\u843C`].string() // U+843C <cjk>
	0xD4: [`\u855A`].string() // U+855A <cjk>
	0xD5: [`\u8484`].string() // U+8484 <cjk>
	0xD6: [`\u8477`].string() // U+8477 <cjk>
	0xD7: [`\u846B`].string() // U+846B <cjk>
	0xD8: [`\u84AD`].string() // U+84AD <cjk>
	0xD9: [`\u846E`].string() // U+846E <cjk>
	0xDA: [`\u8482`].string() // U+8482 <cjk>
	0xDB: [`\u8469`].string() // U+8469 <cjk>
	0xDC: [`\u8446`].string() // U+8446 <cjk>
	0xDD: [`\u842C`].string() // U+842C <cjk>
	0xDE: [`\u846F`].string() // U+846F <cjk>
	0xDF: [`\u8479`].string() // U+8479 <cjk>
	0xE0: [`\u8435`].string() // U+8435 <cjk>
	0xE1: [`\u84CA`].string() // U+84CA <cjk>
	0xE2: [`\u8462`].string() // U+8462 <cjk>
	0xE3: [`\u84B9`].string() // U+84B9 <cjk>
	0xE4: [`\u84BF`].string() // U+84BF <cjk>
	0xE5: [`\u849F`].string() // U+849F <cjk>
	0xE6: [`\u84D9`].string() // U+84D9 <cjk>
	0xE7: [`\u84CD`].string() // U+84CD <cjk>
	0xE8: [`\u84BB`].string() // U+84BB <cjk>
	0xE9: [`\u84DA`].string() // U+84DA <cjk>
	0xEA: [`\u84D0`].string() // U+84D0 <cjk>
	0xEB: [`\u84C1`].string() // U+84C1 <cjk>
	0xEC: [`\u84C6`].string() // U+84C6 <cjk>
	0xED: [`\u84D6`].string() // U+84D6 <cjk>
	0xEE: [`\u84A1`].string() // U+84A1 <cjk>
	0xEF: [`\u8521`].string() // U+8521 <cjk>
	0xF0: [`\u84FF`].string() // U+84FF <cjk>
	0xF1: [`\u84F4`].string() // U+84F4 <cjk>
	0xF2: [`\u8517`].string() // U+8517 <cjk>
	0xF3: [`\u8518`].string() // U+8518 <cjk>
	0xF4: [`\u852C`].string() // U+852C <cjk>
	0xF5: [`\u851F`].string() // U+851F <cjk>
	0xF6: [`\u8515`].string() // U+8515 <cjk>
	0xF7: [`\u8514`].string() // U+8514 <cjk>
	0xF8: [`\u84FC`].string() // U+84FC <cjk>
	0xF9: [`\u8540`].string() // U+8540 <cjk>
	0xFA: [`\u8563`].string() // U+8563 <cjk>
	0xFB: [`\u8558`].string() // U+8558 <cjk>
	0xFC: [`\u8548`].string() // U+8548 <cjk>
}

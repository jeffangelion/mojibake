module mojibake

const jis_x_0213_doublebyte_0x8f = {
	0x40: [`\u5B97`].string() // U+5B97 <cjk>
	0x41: [`\u5C31`].string() // U+5C31 <cjk>
	0x42: [`\u5DDE`].string() // U+5DDE <cjk>
	0x43: [`\u4FEE`].string() // U+4FEE <cjk>
	0x44: [`\u6101`].string() // U+6101 <cjk>
	0x45: [`\u62FE`].string() // U+62FE <cjk>
	0x46: [`\u6D32`].string() // U+6D32 <cjk>
	0x47: [`\u79C0`].string() // U+79C0 <cjk>
	0x48: [`\u79CB`].string() // U+79CB <cjk>
	0x49: [`\u7D42`].string() // U+7D42 <cjk>
	0x4A: [`\u7E4D`].string() // U+7E4D <cjk>
	0x4B: [`\u7FD2`].string() // U+7FD2 <cjk>
	0x4C: [`\u81ED`].string() // U+81ED <cjk>
	0x4D: [`\u821F`].string() // U+821F <cjk>
	0x4E: [`\u8490`].string() // U+8490 <cjk>
	0x4F: [`\u8846`].string() // U+8846 <cjk>
	0x50: [`\u8972`].string() // U+8972 <cjk>
	0x51: [`\u8B90`].string() // U+8B90 <cjk>
	0x52: [`\u8E74`].string() // U+8E74 <cjk>
	0x53: [`\u8F2F`].string() // U+8F2F <cjk>
	0x54: [`\u9031`].string() // U+9031 <cjk>
	0x55: [`\u914B`].string() // U+914B <cjk>
	0x56: [`\u916C`].string() // U+916C <cjk>
	0x57: [`\u96C6`].string() // U+96C6 <cjk>
	0x58: [`\u919C`].string() // U+919C <cjk>
	0x59: [`\u4EC0`].string() // U+4EC0 <cjk>
	0x5A: [`\u4F4F`].string() // U+4F4F <cjk>
	0x5B: [`\u5145`].string() // U+5145 <cjk>
	0x5C: [`\u5341`].string() // U+5341 <cjk>
	0x5D: [`\u5F93`].string() // U+5F93 <cjk>
	0x5E: [`\u620E`].string() // U+620E <cjk>
	0x5F: [`\u67D4`].string() // U+67D4 <cjk>
	0x60: [`\u6C41`].string() // U+6C41 <cjk>
	0x61: [`\u6E0B`].string() // U+6E0B <cjk>
	0x62: [`\u7363`].string() // U+7363 <cjk>
	0x63: [`\u7E26`].string() // U+7E26 <cjk>
	0x64: [`\u91CD`].string() // U+91CD <cjk>
	0x65: [`\u9283`].string() // U+9283 <cjk>
	0x66: [`\u53D4`].string() // U+53D4 <cjk>
	0x67: [`\u5919`].string() // U+5919 <cjk>
	0x68: [`\u5BBF`].string() // U+5BBF <cjk>
	0x69: [`\u6DD1`].string() // U+6DD1 <cjk>
	0x6A: [`\u795D`].string() // U+795D <cjk>
	0x6B: [`\u7E2E`].string() // U+7E2E <cjk>
	0x6C: [`\u7C9B`].string() // U+7C9B <cjk>
	0x6D: [`\u587E`].string() // U+587E <cjk>
	0x6E: [`\u719F`].string() // U+719F <cjk>
	0x6F: [`\u51FA`].string() // U+51FA <cjk>
	0x70: [`\u8853`].string() // U+8853 <cjk>
	0x71: [`\u8FF0`].string() // U+8FF0 <cjk>
	0x72: [`\u4FCA`].string() // U+4FCA <cjk>
	0x73: [`\u5CFB`].string() // U+5CFB <cjk>
	0x74: [`\u6625`].string() // U+6625 <cjk>
	0x75: [`\u77AC`].string() // U+77AC <cjk>
	0x76: [`\u7AE3`].string() // U+7AE3 <cjk>
	0x77: [`\u821C`].string() // U+821C <cjk>
	0x78: [`\u99FF`].string() // U+99FF <cjk>
	0x79: [`\u51C6`].string() // U+51C6 <cjk>
	0x7A: [`\u5FAA`].string() // U+5FAA <cjk>
	0x7B: [`\u65EC`].string() // U+65EC <cjk>
	0x7C: [`\u696F`].string() // U+696F <cjk>
	0x7D: [`\u6B89`].string() // U+6B89 <cjk>
	0x7E: [`\u6DF3`].string() // U+6DF3 <cjk>
	0x80: [`\u6E96`].string() // U+6E96 <cjk>
	0x81: [`\u6F64`].string() // U+6F64 <cjk>
	0x82: [`\u76FE`].string() // U+76FE <cjk>
	0x83: [`\u7D14`].string() // U+7D14 <cjk>
	0x84: [`\u5DE1`].string() // U+5DE1 <cjk>
	0x85: [`\u9075`].string() // U+9075 <cjk>
	0x86: [`\u9187`].string() // U+9187 <cjk>
	0x87: [`\u9806`].string() // U+9806 <cjk>
	0x88: [`\u51E6`].string() // U+51E6 <cjk>
	0x89: [`\u521D`].string() // U+521D <cjk>
	0x8A: [`\u6240`].string() // U+6240 <cjk>
	0x8B: [`\u6691`].string() // U+6691 <cjk>
	0x8C: [`\u66D9`].string() // U+66D9 <cjk>
	0x8D: [`\u6E1A`].string() // U+6E1A <cjk>
	0x8E: [`\u5EB6`].string() // U+5EB6 <cjk>
	0x8F: [`\u7DD2`].string() // U+7DD2 <cjk>
	0x90: [`\u7F72`].string() // U+7F72 <cjk>
	0x91: [`\u66F8`].string() // U+66F8 <cjk>
	0x92: [`\u85AF`].string() // U+85AF <cjk>
	0x93: [`\u85F7`].string() // U+85F7 <cjk>
	0x94: [`\u8AF8`].string() // U+8AF8 <cjk>
	0x95: [`\u52A9`].string() // U+52A9 <cjk>
	0x96: [`\u53D9`].string() // U+53D9 <cjk>
	0x97: [`\u5973`].string() // U+5973 <cjk>
	0x98: [`\u5E8F`].string() // U+5E8F <cjk>
	0x99: [`\u5F90`].string() // U+5F90 <cjk>
	0x9A: [`\u6055`].string() // U+6055 <cjk>
	0x9B: [`\u92E4`].string() // U+92E4 <cjk>
	0x9C: [`\u9664`].string() // U+9664 <cjk>
	0x9D: [`\u50B7`].string() // U+50B7 <cjk>
	0x9E: [`\u511F`].string() // U+511F <cjk>
	0x9F: [`\u52DD`].string() // U+52DD <cjk>
	0xA0: [`\u5320`].string() // U+5320 <cjk>
	0xA1: [`\u5347`].string() // U+5347 <cjk>
	0xA2: [`\u53EC`].string() // U+53EC <cjk>
	0xA3: [`\u54E8`].string() // U+54E8 <cjk>
	0xA4: [`\u5546`].string() // U+5546 <cjk>
	0xA5: [`\u5531`].string() // U+5531 <cjk>
	0xA6: [`\u5617`].string() // U+5617 <cjk>
	0xA7: [`\u5968`].string() // U+5968 <cjk>
	0xA8: [`\u59BE`].string() // U+59BE <cjk>
	0xA9: [`\u5A3C`].string() // U+5A3C <cjk>
	0xAA: [`\u5BB5`].string() // U+5BB5 <cjk>
	0xAB: [`\u5C06`].string() // U+5C06 <cjk>
	0xAC: [`\u5C0F`].string() // U+5C0F <cjk>
	0xAD: [`\u5C11`].string() // U+5C11 <cjk>
	0xAE: [`\u5C1A`].string() // U+5C1A <cjk>
	0xAF: [`\u5E84`].string() // U+5E84 <cjk>
	0xB0: [`\u5E8A`].string() // U+5E8A <cjk>
	0xB1: [`\u5EE0`].string() // U+5EE0 <cjk>
	0xB2: [`\u5F70`].string() // U+5F70 <cjk>
	0xB3: [`\u627F`].string() // U+627F <cjk>
	0xB4: [`\u6284`].string() // U+6284 <cjk>
	0xB5: [`\u62DB`].string() // U+62DB <cjk>
	0xB6: [`\u638C`].string() // U+638C <cjk>
	0xB7: [`\u6377`].string() // U+6377 <cjk>
	0xB8: [`\u6607`].string() // U+6607 <cjk>
	0xB9: [`\u660C`].string() // U+660C <cjk>
	0xBA: [`\u662D`].string() // U+662D <cjk>
	0xBB: [`\u6676`].string() // U+6676 <cjk>
	0xBC: [`\u677E`].string() // U+677E <cjk>
	0xBD: [`\u68A2`].string() // U+68A2 <cjk>
	0xBE: [`\u6A1F`].string() // U+6A1F <cjk>
	0xBF: [`\u6A35`].string() // U+6A35 <cjk>
	0xC0: [`\u6CBC`].string() // U+6CBC <cjk>
	0xC1: [`\u6D88`].string() // U+6D88 <cjk>
	0xC2: [`\u6E09`].string() // U+6E09 <cjk>
	0xC3: [`\u6E58`].string() // U+6E58 <cjk>
	0xC4: [`\u713C`].string() // U+713C <cjk>
	0xC5: [`\u7126`].string() // U+7126 <cjk>
	0xC6: [`\u7167`].string() // U+7167 <cjk>
	0xC7: [`\u75C7`].string() // U+75C7 <cjk>
	0xC8: [`\u7701`].string() // U+7701 <cjk>
	0xC9: [`\u785D`].string() // U+785D <cjk>
	0xCA: [`\u7901`].string() // U+7901 <cjk>
	0xCB: [`\u7965`].string() // U+7965 <cjk>
	0xCC: [`\u79F0`].string() // U+79F0 <cjk>
	0xCD: [`\u7AE0`].string() // U+7AE0 <cjk>
	0xCE: [`\u7B11`].string() // U+7B11 <cjk>
	0xCF: [`\u7CA7`].string() // U+7CA7 <cjk>
	0xD0: [`\u7D39`].string() // U+7D39 <cjk>
	0xD1: [`\u8096`].string() // U+8096 <cjk>
	0xD2: [`\u83D6`].string() // U+83D6 <cjk>
	0xD3: [`\u848B`].string() // U+848B <cjk>
	0xD4: [`\u8549`].string() // U+8549 <cjk>
	0xD5: [`\u885D`].string() // U+885D <cjk>
	0xD6: [`\u88F3`].string() // U+88F3 <cjk>
	0xD7: [`\u8A1F`].string() // U+8A1F <cjk>
	0xD8: [`\u8A3C`].string() // U+8A3C <cjk>
	0xD9: [`\u8A54`].string() // U+8A54 <cjk>
	0xDA: [`\u8A73`].string() // U+8A73 <cjk>
	0xDB: [`\u8C61`].string() // U+8C61 <cjk>
	0xDC: [`\u8CDE`].string() // U+8CDE <cjk>
	0xDD: [`\u91A4`].string() // U+91A4 <cjk>
	0xDE: [`\u9266`].string() // U+9266 <cjk>
	0xDF: [`\u937E`].string() // U+937E <cjk>
	0xE0: [`\u9418`].string() // U+9418 <cjk>
	0xE1: [`\u969C`].string() // U+969C <cjk>
	0xE2: [`\u9798`].string() // U+9798 <cjk>
	0xE3: [`\u4E0A`].string() // U+4E0A <cjk>
	0xE4: [`\u4E08`].string() // U+4E08 <cjk>
	0xE5: [`\u4E1E`].string() // U+4E1E <cjk>
	0xE6: [`\u4E57`].string() // U+4E57 <cjk>
	0xE7: [`\u5197`].string() // U+5197 <cjk>
	0xE8: [`\u5270`].string() // U+5270 <cjk>
	0xE9: [`\u57CE`].string() // U+57CE <cjk>
	0xEA: [`\u5834`].string() // U+5834 <cjk>
	0xEB: [`\u58CC`].string() // U+58CC <cjk>
	0xEC: [`\u5B22`].string() // U+5B22 <cjk>
	0xED: [`\u5E38`].string() // U+5E38 <cjk>
	0xEE: [`\u60C5`].string() // U+60C5 <cjk>
	0xEF: [`\u64FE`].string() // U+64FE <cjk>
	0xF0: [`\u6761`].string() // U+6761 <cjk>
	0xF1: [`\u6756`].string() // U+6756 <cjk>
	0xF2: [`\u6D44`].string() // U+6D44 <cjk>
	0xF3: [`\u72B6`].string() // U+72B6 <cjk>
	0xF4: [`\u7573`].string() // U+7573 <cjk>
	0xF5: [`\u7A63`].string() // U+7A63 <cjk>
	0xF6: [`\u84B8`].string() // U+84B8 <cjk>
	0xF7: [`\u8B72`].string() // U+8B72 <cjk>
	0xF8: [`\u91B8`].string() // U+91B8 <cjk>
	0xF9: [`\u9320`].string() // U+9320 <cjk>
	0xFA: [`\u5631`].string() // U+5631 <cjk>
	0xFB: [`\u57F4`].string() // U+57F4 <cjk>
	0xFC: [`\u98FE`].string() // U+98FE <cjk>
}

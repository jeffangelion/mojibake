module mojibake

const jis_x_0213_doublebyte_0x91 = {
	0x40: [`\u7E4A`].string() // U+7E4A <cjk>
	0x41: [`\u7FA8`].string() // U+7FA8 <cjk>
	0x42: [`\u817A`].string() // U+817A <cjk>
	0x43: [`\u821B`].string() // U+821B <cjk>
	0x44: [`\u8239`].string() // U+8239 <cjk>
	0x45: [`\u85A6`].string() // U+85A6 <cjk>
	0x46: [`\u8A6E`].string() // U+8A6E <cjk>
	0x47: [`\u8CCE`].string() // U+8CCE <cjk>
	0x48: [`\u8DF5`].string() // U+8DF5 <cjk>
	0x49: [`\u9078`].string() // U+9078 <cjk>
	0x4A: [`\u9077`].string() // U+9077 <cjk>
	0x4B: [`\u92AD`].string() // U+92AD <cjk>
	0x4C: [`\u9291`].string() // U+9291 <cjk>
	0x4D: [`\u9583`].string() // U+9583 <cjk>
	0x4E: [`\u9BAE`].string() // U+9BAE <cjk>
	0x4F: [`\u524D`].string() // U+524D <cjk>
	0x50: [`\u5584`].string() // U+5584 <cjk>
	0x51: [`\u6F38`].string() // U+6F38 <cjk>
	0x52: [`\u7136`].string() // U+7136 <cjk>
	0x53: [`\u5168`].string() // U+5168 <cjk>
	0x54: [`\u7985`].string() // U+7985 <cjk>
	0x55: [`\u7E55`].string() // U+7E55 <cjk>
	0x56: [`\u81B3`].string() // U+81B3 <cjk>
	0x57: [`\u7CCE`].string() // U+7CCE <cjk>
	0x58: [`\u564C`].string() // U+564C <cjk>
	0x59: [`\u5851`].string() // U+5851 <cjk>
	0x5A: [`\u5CA8`].string() // U+5CA8 <cjk>
	0x5B: [`\u63AA`].string() // U+63AA <cjk>
	0x5C: [`\u66FE`].string() // U+66FE <cjk>
	0x5D: [`\u66FD`].string() // U+66FD <cjk>
	0x5E: [`\u695A`].string() // U+695A <cjk>
	0x5F: [`\u72D9`].string() // U+72D9 <cjk>
	0x60: [`\u758F`].string() // U+758F <cjk>
	0x61: [`\u758E`].string() // U+758E <cjk>
	0x62: [`\u790E`].string() // U+790E <cjk>
	0x63: [`\u7956`].string() // U+7956 <cjk>
	0x64: [`\u79DF`].string() // U+79DF <cjk>
	0x65: [`\u7C97`].string() // U+7C97 <cjk>
	0x66: [`\u7D20`].string() // U+7D20 <cjk>
	0x67: [`\u7D44`].string() // U+7D44 <cjk>
	0x68: [`\u8607`].string() // U+8607 <cjk>
	0x69: [`\u8A34`].string() // U+8A34 <cjk>
	0x6A: [`\u963B`].string() // U+963B <cjk>
	0x6B: [`\u9061`].string() // U+9061 <cjk>
	0x6C: [`\u9F20`].string() // U+9F20 <cjk>
	0x6D: [`\u50E7`].string() // U+50E7 <cjk>
	0x6E: [`\u5275`].string() // U+5275 <cjk>
	0x6F: [`\u53CC`].string() // U+53CC <cjk>
	0x70: [`\u53E2`].string() // U+53E2 <cjk>
	0x71: [`\u5009`].string() // U+5009 <cjk>
	0x72: [`\u55AA`].string() // U+55AA <cjk>
	0x73: [`\u58EE`].string() // U+58EE <cjk>
	0x74: [`\u594F`].string() // U+594F <cjk>
	0x75: [`\u723D`].string() // U+723D <cjk>
	0x76: [`\u5B8B`].string() // U+5B8B <cjk>
	0x77: [`\u5C64`].string() // U+5C64 <cjk>
	0x78: [`\u531D`].string() // U+531D <cjk>
	0x79: [`\u60E3`].string() // U+60E3 <cjk>
	0x7A: [`\u60F3`].string() // U+60F3 <cjk>
	0x7B: [`\u635C`].string() // U+635C <cjk>
	0x7C: [`\u6383`].string() // U+6383 <cjk>
	0x7D: [`\u633F`].string() // U+633F <cjk>
	0x7E: [`\u63BB`].string() // U+63BB <cjk>
	0x80: [`\u64CD`].string() // U+64CD <cjk>
	0x81: [`\u65E9`].string() // U+65E9 <cjk>
	0x82: [`\u66F9`].string() // U+66F9 <cjk>
	0x83: [`\u5DE3`].string() // U+5DE3 <cjk>
	0x84: [`\u69CD`].string() // U+69CD <cjk>
	0x85: [`\u69FD`].string() // U+69FD <cjk>
	0x86: [`\u6F15`].string() // U+6F15 <cjk>
	0x87: [`\u71E5`].string() // U+71E5 <cjk>
	0x88: [`\u4E89`].string() // U+4E89 <cjk>
	0x89: [`\u75E9`].string() // U+75E9 <cjk>
	0x8A: [`\u76F8`].string() // U+76F8 <cjk>
	0x8B: [`\u7A93`].string() // U+7A93 <cjk>
	0x8C: [`\u7CDF`].string() // U+7CDF <cjk>
	0x8D: [`\u7DCF`].string() // U+7DCF <cjk>
	0x8E: [`\u7D9C`].string() // U+7D9C <cjk>
	0x8F: [`\u8061`].string() // U+8061 <cjk>
	0x90: [`\u8349`].string() // U+8349 <cjk>
	0x91: [`\u8358`].string() // U+8358 <cjk>
	0x92: [`\u846C`].string() // U+846C <cjk>
	0x93: [`\u84BC`].string() // U+84BC <cjk>
	0x94: [`\u85FB`].string() // U+85FB <cjk>
	0x95: [`\u88C5`].string() // U+88C5 <cjk>
	0x96: [`\u8D70`].string() // U+8D70 <cjk>
	0x97: [`\u9001`].string() // U+9001 <cjk>
	0x98: [`\u906D`].string() // U+906D <cjk>
	0x99: [`\u9397`].string() // U+9397 <cjk>
	0x9A: [`\u971C`].string() // U+971C <cjk>
	0x9B: [`\u9A12`].string() // U+9A12 <cjk>
	0x9C: [`\u50CF`].string() // U+50CF <cjk>
	0x9D: [`\u5897`].string() // U+5897 <cjk>
	0x9E: [`\u618E`].string() // U+618E <cjk>
	0x9F: [`\u81D3`].string() // U+81D3 <cjk>
	0xA0: [`\u8535`].string() // U+8535 <cjk>
	0xA1: [`\u8D08`].string() // U+8D08 <cjk>
	0xA2: [`\u9020`].string() // U+9020 <cjk>
	0xA3: [`\u4FC3`].string() // U+4FC3 <cjk>
	0xA4: [`\u5074`].string() // U+5074 <cjk>
	0xA5: [`\u5247`].string() // U+5247 <cjk>
	0xA6: [`\u5373`].string() // U+5373 <cjk>
	0xA7: [`\u606F`].string() // U+606F <cjk>
	0xA8: [`\u6349`].string() // U+6349 <cjk>
	0xA9: [`\u675F`].string() // U+675F <cjk>
	0xAA: [`\u6E2C`].string() // U+6E2C <cjk>
	0xAB: [`\u8DB3`].string() // U+8DB3 <cjk>
	0xAC: [`\u901F`].string() // U+901F <cjk>
	0xAD: [`\u4FD7`].string() // U+4FD7 <cjk>
	0xAE: [`\u5C5E`].string() // U+5C5E <cjk>
	0xAF: [`\u8CCA`].string() // U+8CCA <cjk>
	0xB0: [`\u65CF`].string() // U+65CF <cjk>
	0xB1: [`\u7D9A`].string() // U+7D9A <cjk>
	0xB2: [`\u5352`].string() // U+5352 <cjk>
	0xB3: [`\u8896`].string() // U+8896 <cjk>
	0xB4: [`\u5176`].string() // U+5176 <cjk>
	0xB5: [`\u63C3`].string() // U+63C3 <cjk>
	0xB6: [`\u5B58`].string() // U+5B58 <cjk>
	0xB7: [`\u5B6B`].string() // U+5B6B <cjk>
	0xB8: [`\u5C0A`].string() // U+5C0A <cjk>
	0xB9: [`\u640D`].string() // U+640D <cjk>
	0xBA: [`\u6751`].string() // U+6751 <cjk>
	0xBB: [`\u905C`].string() // U+905C <cjk>
	0xBC: [`\u4ED6`].string() // U+4ED6 <cjk>
	0xBD: [`\u591A`].string() // U+591A <cjk>
	0xBE: [`\u592A`].string() // U+592A <cjk>
	0xBF: [`\u6C70`].string() // U+6C70 <cjk>
	0xC0: [`\u8A51`].string() // U+8A51 <cjk>
	0xC1: [`\u553E`].string() // U+553E <cjk>
	0xC2: [`\u5815`].string() // U+5815 <cjk>
	0xC3: [`\u59A5`].string() // U+59A5 <cjk>
	0xC4: [`\u60F0`].string() // U+60F0 <cjk>
	0xC5: [`\u6253`].string() // U+6253 <cjk>
	0xC6: [`\u67C1`].string() // U+67C1 <cjk>
	0xC7: [`\u8235`].string() // U+8235 <cjk>
	0xC8: [`\u6955`].string() // U+6955 <cjk>
	0xC9: [`\u9640`].string() // U+9640 <cjk>
	0xCA: [`\u99C4`].string() // U+99C4 <cjk>
	0xCB: [`\u9A28`].string() // U+9A28 <cjk>
	0xCC: [`\u4F53`].string() // U+4F53 <cjk>
	0xCD: [`\u5806`].string() // U+5806 <cjk>
	0xCE: [`\u5BFE`].string() // U+5BFE <cjk>
	0xCF: [`\u8010`].string() // U+8010 <cjk>
	0xD0: [`\u5CB1`].string() // U+5CB1 <cjk>
	0xD1: [`\u5E2F`].string() // U+5E2F <cjk>
	0xD2: [`\u5F85`].string() // U+5F85 <cjk>
	0xD3: [`\u6020`].string() // U+6020 <cjk>
	0xD4: [`\u614B`].string() // U+614B <cjk>
	0xD5: [`\u6234`].string() // U+6234 <cjk>
	0xD6: [`\u66FF`].string() // U+66FF <cjk>
	0xD7: [`\u6CF0`].string() // U+6CF0 <cjk>
	0xD8: [`\u6EDE`].string() // U+6EDE <cjk>
	0xD9: [`\u80CE`].string() // U+80CE <cjk>
	0xDA: [`\u817F`].string() // U+817F <cjk>
	0xDB: [`\u82D4`].string() // U+82D4 <cjk>
	0xDC: [`\u888B`].string() // U+888B <cjk>
	0xDD: [`\u8CB8`].string() // U+8CB8 <cjk>
	0xDE: [`\u9000`].string() // U+9000 <cjk>
	0xDF: [`\u902E`].string() // U+902E <cjk>
	0xE0: [`\u968A`].string() // U+968A <cjk>
	0xE1: [`\u9EDB`].string() // U+9EDB <cjk>
	0xE2: [`\u9BDB`].string() // U+9BDB <cjk>
	0xE3: [`\u4EE3`].string() // U+4EE3 <cjk>
	0xE4: [`\u53F0`].string() // U+53F0 <cjk>
	0xE5: [`\u5927`].string() // U+5927 <cjk>
	0xE6: [`\u7B2C`].string() // U+7B2C <cjk>
	0xE7: [`\u918D`].string() // U+918D <cjk>
	0xE8: [`\u984C`].string() // U+984C <cjk>
	0xE9: [`\u9DF9`].string() // U+9DF9 <cjk>
	0xEA: [`\u6EDD`].string() // U+6EDD <cjk>
	0xEB: [`\u7027`].string() // U+7027 <cjk>
	0xEC: [`\u5353`].string() // U+5353 <cjk>
	0xED: [`\u5544`].string() // U+5544 <cjk>
	0xEE: [`\u5B85`].string() // U+5B85 <cjk>
	0xEF: [`\u6258`].string() // U+6258 <cjk>
	0xF0: [`\u629E`].string() // U+629E <cjk>
	0xF1: [`\u62D3`].string() // U+62D3 <cjk>
	0xF2: [`\u6CA2`].string() // U+6CA2 <cjk>
	0xF3: [`\u6FEF`].string() // U+6FEF <cjk>
	0xF4: [`\u7422`].string() // U+7422 <cjk>
	0xF5: [`\u8A17`].string() // U+8A17 <cjk>
	0xF6: [`\u9438`].string() // U+9438 <cjk>
	0xF7: [`\u6FC1`].string() // U+6FC1 <cjk>
	0xF8: [`\u8AFE`].string() // U+8AFE <cjk>
	0xF9: [`\u8338`].string() // U+8338 <cjk>
	0xFA: [`\u51E7`].string() // U+51E7 <cjk>
	0xFB: [`\u86F8`].string() // U+86F8 <cjk>
	0xFC: [`\u53EA`].string() // U+53EA <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xf0 = {
	0x40: utf32_to_str(0x20089) // U+20089 <cjk>
	0x41: [`\u4E02`].string() // U+4E02 <cjk>
	0x42: [`\u4E0F`].string() // U+4E0F <cjk>
	0x43: [`\u4E12`].string() // U+4E12 <cjk>
	0x44: [`\u4E29`].string() // U+4E29 <cjk>
	0x45: [`\u4E2B`].string() // U+4E2B <cjk>
	0x46: [`\u4E2E`].string() // U+4E2E <cjk>
	0x47: [`\u4E40`].string() // U+4E40 <cjk>
	0x48: [`\u4E47`].string() // U+4E47 <cjk>
	0x49: [`\u4E48`].string() // U+4E48 <cjk>
	0x4A: utf32_to_str(0x200A2) // U+200A2 <cjk>
	0x4B: [`\u4E51`].string() // U+4E51 <cjk>
	0x4C: [`\u3406`].string() // U+3406 <cjk>
	0x4D: utf32_to_str(0x200A4) // U+200A4 <cjk>
	0x4E: [`\u4E5A`].string() // U+4E5A <cjk>
	0x4F: [`\u4E69`].string() // U+4E69 <cjk>
	0x50: [`\u4E9D`].string() // U+4E9D <cjk>
	0x51: [`\u342C`].string() // U+342C <cjk>
	0x52: [`\u342E`].string() // U+342E <cjk>
	0x53: [`\u4EB9`].string() // U+4EB9 <cjk>
	0x54: [`\u4EBB`].string() // U+4EBB <cjk>
	0x55: utf32_to_str(0x201A2) // U+201A2 <cjk>
	0x56: [`\u4EBC`].string() // U+4EBC <cjk>
	0x57: [`\u4EC3`].string() // U+4EC3 <cjk>
	0x58: [`\u4EC8`].string() // U+4EC8 <cjk>
	0x59: [`\u4ED0`].string() // U+4ED0 <cjk>
	0x5A: [`\u4EEB`].string() // U+4EEB <cjk>
	0x5B: [`\u4EDA`].string() // U+4EDA <cjk>
	0x5C: [`\u4EF1`].string() // U+4EF1 <cjk>
	0x5D: [`\u4EF5`].string() // U+4EF5 <cjk>
	0x5E: [`\u4F00`].string() // U+4F00 <cjk>
	0x5F: [`\u4F16`].string() // U+4F16 <cjk>
	0x60: [`\u4F64`].string() // U+4F64 <cjk>
	0x61: [`\u4F37`].string() // U+4F37 <cjk>
	0x62: [`\u4F3E`].string() // U+4F3E <cjk>
	0x63: [`\u4F54`].string() // U+4F54 <cjk>
	0x64: [`\u4F58`].string() // U+4F58 <cjk>
	0x65: utf32_to_str(0x20213) // U+20213 <cjk>
	0x66: [`\u4F77`].string() // U+4F77 <cjk>
	0x67: [`\u4F78`].string() // U+4F78 <cjk>
	0x68: [`\u4F7A`].string() // U+4F7A <cjk>
	0x69: [`\u4F7D`].string() // U+4F7D <cjk>
	0x6A: [`\u4F82`].string() // U+4F82 <cjk>
	0x6B: [`\u4F85`].string() // U+4F85 <cjk>
	0x6C: [`\u4F92`].string() // U+4F92 <cjk>
	0x6D: [`\u4F9A`].string() // U+4F9A <cjk>
	0x6E: [`\u4FE6`].string() // U+4FE6 <cjk>
	0x6F: [`\u4FB2`].string() // U+4FB2 <cjk>
	0x70: [`\u4FBE`].string() // U+4FBE <cjk>
	0x71: [`\u4FC5`].string() // U+4FC5 <cjk>
	0x72: [`\u4FCB`].string() // U+4FCB <cjk>
	0x73: [`\u4FCF`].string() // U+4FCF <cjk>
	0x74: [`\u4FD2`].string() // U+4FD2 <cjk>
	0x75: [`\u346A`].string() // U+346A <cjk>
	0x76: [`\u4FF2`].string() // U+4FF2 <cjk>
	0x77: [`\u5000`].string() // U+5000 <cjk>
	0x78: [`\u5010`].string() // U+5010 <cjk>
	0x79: [`\u5013`].string() // U+5013 <cjk>
	0x7A: [`\u501C`].string() // U+501C <cjk>
	0x7B: [`\u501E`].string() // U+501E <cjk>
	0x7C: [`\u5022`].string() // U+5022 <cjk>
	0x7D: [`\u3468`].string() // U+3468 <cjk>
	0x7E: [`\u5042`].string() // U+5042 <cjk>
	0x80: [`\u5046`].string() // U+5046 <cjk>
	0x81: [`\u504E`].string() // U+504E <cjk>
	0x82: [`\u5053`].string() // U+5053 <cjk>
	0x83: [`\u5057`].string() // U+5057 <cjk>
	0x84: [`\u5063`].string() // U+5063 <cjk>
	0x85: [`\u5066`].string() // U+5066 <cjk>
	0x86: [`\u506A`].string() // U+506A <cjk>
	0x87: [`\u5070`].string() // U+5070 <cjk>
	0x88: [`\u50A3`].string() // U+50A3 <cjk>
	0x89: [`\u5088`].string() // U+5088 <cjk>
	0x8A: [`\u5092`].string() // U+5092 <cjk>
	0x8B: [`\u5093`].string() // U+5093 <cjk>
	0x8C: [`\u5095`].string() // U+5095 <cjk>
	0x8D: [`\u5096`].string() // U+5096 <cjk>
	0x8E: [`\u509C`].string() // U+509C <cjk>
	0x8F: [`\u50AA`].string() // U+50AA <cjk>
	0x90: utf32_to_str(0x2032B) // U+2032B <cjk>
	0x91: [`\u50B1`].string() // U+50B1 <cjk>
	0x92: [`\u50BA`].string() // U+50BA <cjk>
	0x93: [`\u50BB`].string() // U+50BB <cjk>
	0x94: [`\u50C4`].string() // U+50C4 <cjk>
	0x95: [`\u50C7`].string() // U+50C7 <cjk>
	0x96: [`\u50F3`].string() // U+50F3 <cjk>
	0x97: utf32_to_str(0x20381) // U+20381 <cjk>
	0x98: [`\u50CE`].string() // U+50CE <cjk>
	0x99: utf32_to_str(0x20371) // U+20371 <cjk>
	0x9A: [`\u50D4`].string() // U+50D4 <cjk>
	0x9B: [`\u50D9`].string() // U+50D9 <cjk>
	0x9C: [`\u50E1`].string() // U+50E1 <cjk>
	0x9D: [`\u50E9`].string() // U+50E9 <cjk>
	0x9E: [`\u3492`].string() // U+3492 <cjk>
	0x9F: [`\u5B96`].string() // U+5B96 <cjk>
	0xA0: [`\u5BAC`].string() // U+5BAC <cjk>
	0xA1: [`\u3761`].string() // U+3761 <cjk>
	0xA2: [`\u5BC0`].string() // U+5BC0 <cjk>
	0xA3: [`\u3762`].string() // U+3762 <cjk>
	0xA4: [`\u5BCE`].string() // U+5BCE <cjk>
	0xA5: [`\u5BD6`].string() // U+5BD6 <cjk>
	0xA6: [`\u376C`].string() // U+376C <cjk>
	0xA7: [`\u376B`].string() // U+376B <cjk>
	0xA8: [`\u5BF1`].string() // U+5BF1 <cjk>
	0xA9: [`\u5BFD`].string() // U+5BFD <cjk>
	0xAA: [`\u3775`].string() // U+3775 <cjk>
	0xAB: [`\u5C03`].string() // U+5C03 <cjk>
	0xAC: [`\u5C29`].string() // U+5C29 <cjk>
	0xAD: [`\u5C30`].string() // U+5C30 <cjk>
	0xAE: utf32_to_str(0x21C56) // U+21C56 <cjk>
	0xAF: [`\u5C5F`].string() // U+5C5F <cjk>
	0xB0: [`\u5C63`].string() // U+5C63 <cjk>
	0xB1: [`\u5C67`].string() // U+5C67 <cjk>
	0xB2: [`\u5C68`].string() // U+5C68 <cjk>
	0xB3: [`\u5C69`].string() // U+5C69 <cjk>
	0xB4: [`\u5C70`].string() // U+5C70 <cjk>
	0xB5: utf32_to_str(0x21D2D) // U+21D2D <cjk>
	0xB6: utf32_to_str(0x21D45) // U+21D45 <cjk>
	0xB7: [`\u5C7C`].string() // U+5C7C <cjk>
	0xB8: utf32_to_str(0x21D78) // U+21D78 <cjk>
	0xB9: utf32_to_str(0x21D62) // U+21D62 <cjk>
	0xBA: [`\u5C88`].string() // U+5C88 <cjk>
	0xBB: [`\u5C8A`].string() // U+5C8A <cjk>
	0xBC: [`\u37C1`].string() // U+37C1 <cjk>
	0xBD: utf32_to_str(0x21DA1) // U+21DA1 <cjk>
	0xBE: utf32_to_str(0x21D9C) // U+21D9C <cjk>
	0xBF: [`\u5CA0`].string() // U+5CA0 <cjk>
	0xC0: [`\u5CA2`].string() // U+5CA2 <cjk>
	0xC1: [`\u5CA6`].string() // U+5CA6 <cjk>
	0xC2: [`\u5CA7`].string() // U+5CA7 <cjk>
	0xC3: utf32_to_str(0x21D92) // U+21D92 <cjk>
	0xC4: [`\u5CAD`].string() // U+5CAD <cjk>
	0xC5: [`\u5CB5`].string() // U+5CB5 <cjk>
	0xC6: utf32_to_str(0x21DB7) // U+21DB7 <cjk>
	0xC7: [`\u5CC9`].string() // U+5CC9 <cjk>
	0xC8: utf32_to_str(0x21DE0) // U+21DE0 <cjk>
	0xC9: utf32_to_str(0x21E33) // U+21E33 <cjk>
	0xCA: [`\u5D06`].string() // U+5D06 <cjk>
	0xCB: [`\u5D10`].string() // U+5D10 <cjk>
	0xCC: [`\u5D2B`].string() // U+5D2B <cjk>
	0xCD: [`\u5D1D`].string() // U+5D1D <cjk>
	0xCE: [`\u5D20`].string() // U+5D20 <cjk>
	0xCF: [`\u5D24`].string() // U+5D24 <cjk>
	0xD0: [`\u5D26`].string() // U+5D26 <cjk>
	0xD1: [`\u5D31`].string() // U+5D31 <cjk>
	0xD2: [`\u5D39`].string() // U+5D39 <cjk>
	0xD3: [`\u5D42`].string() // U+5D42 <cjk>
	0xD4: [`\u37E8`].string() // U+37E8 <cjk>
	0xD5: [`\u5D61`].string() // U+5D61 <cjk>
	0xD6: [`\u5D6A`].string() // U+5D6A <cjk>
	0xD7: [`\u37F4`].string() // U+37F4 <cjk>
	0xD8: [`\u5D70`].string() // U+5D70 <cjk>
	0xD9: utf32_to_str(0x21F1E) // U+21F1E <cjk>
	0xDA: [`\u37FD`].string() // U+37FD <cjk>
	0xDB: [`\u5D88`].string() // U+5D88 <cjk>
	0xDC: [`\u3800`].string() // U+3800 <cjk>
	0xDD: [`\u5D92`].string() // U+5D92 <cjk>
	0xDE: [`\u5D94`].string() // U+5D94 <cjk>
	0xDF: [`\u5D97`].string() // U+5D97 <cjk>
	0xE0: [`\u5D99`].string() // U+5D99 <cjk>
	0xE1: [`\u5DB0`].string() // U+5DB0 <cjk>
	0xE2: [`\u5DB2`].string() // U+5DB2 <cjk>
	0xE3: [`\u5DB4`].string() // U+5DB4 <cjk>
	0xE4: utf32_to_str(0x21F76) // U+21F76 <cjk>
	0xE5: [`\u5DB9`].string() // U+5DB9 <cjk>
	0xE6: [`\u5DD1`].string() // U+5DD1 <cjk>
	0xE7: [`\u5DD7`].string() // U+5DD7 <cjk>
	0xE8: [`\u5DD8`].string() // U+5DD8 <cjk>
	0xE9: [`\u5DE0`].string() // U+5DE0 <cjk>
	0xEA: utf32_to_str(0x21FFA) // U+21FFA <cjk>
	0xEB: [`\u5DE4`].string() // U+5DE4 <cjk>
	0xEC: [`\u5DE9`].string() // U+5DE9 <cjk>
	0xED: [`\u382F`].string() // U+382F <cjk>
	0xEE: [`\u5E00`].string() // U+5E00 <cjk>
	0xEF: [`\u3836`].string() // U+3836 <cjk>
	0xF0: [`\u5E12`].string() // U+5E12 <cjk>
	0xF1: [`\u5E15`].string() // U+5E15 <cjk>
	0xF2: [`\u3840`].string() // U+3840 <cjk>
	0xF3: [`\u5E1F`].string() // U+5E1F <cjk>
	0xF4: [`\u5E2E`].string() // U+5E2E <cjk>
	0xF5: [`\u5E3E`].string() // U+5E3E <cjk>
	0xF6: [`\u5E49`].string() // U+5E49 <cjk>
	0xF7: [`\u385C`].string() // U+385C <cjk>
	0xF8: [`\u5E56`].string() // U+5E56 <cjk>
	0xF9: [`\u3861`].string() // U+3861 <cjk>
	0xFA: [`\u5E6B`].string() // U+5E6B <cjk>
	0xFB: [`\u5E6C`].string() // U+5E6C <cjk>
	0xFC: [`\u5E6D`].string() // U+5E6D <cjk>
}

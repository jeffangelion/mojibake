module mojibake

const jis_x_0213_doublebyte_0xf3 = {
	0x40: [`\u6299`].string() // U+6299 <cjk>
	0x41: [`\u62A6`].string() // U+62A6 <cjk>
	0x42: [`\u62D5`].string() // U+62D5 <cjk>
	0x43: utf32_to_str(0x22AB8) // U+22AB8 <cjk>
	0x44: [`\u62FD`].string() // U+62FD <cjk>
	0x45: [`\u6303`].string() // U+6303 <cjk>
	0x46: [`\u630D`].string() // U+630D <cjk>
	0x47: [`\u6310`].string() // U+6310 <cjk>
	0x48: utf32_to_str(0x22B4F) // U+22B4F <cjk>
	0x49: utf32_to_str(0x22B50) // U+22B50 <cjk>
	0x4A: [`\u6332`].string() // U+6332 <cjk>
	0x4B: [`\u6335`].string() // U+6335 <cjk>
	0x4C: [`\u633B`].string() // U+633B <cjk>
	0x4D: [`\u633C`].string() // U+633C <cjk>
	0x4E: [`\u6341`].string() // U+6341 <cjk>
	0x4F: [`\u6344`].string() // U+6344 <cjk>
	0x50: [`\u634E`].string() // U+634E <cjk>
	0x51: utf32_to_str(0x22B46) // U+22B46 <cjk>
	0x52: [`\u6359`].string() // U+6359 <cjk>
	0x53: utf32_to_str(0x22C1D) // U+22C1D <cjk>
	0x54: utf32_to_str(0x22BA6) // U+22BA6 <cjk>
	0x55: [`\u636C`].string() // U+636C <cjk>
	0x56: [`\u6384`].string() // U+6384 <cjk>
	0x57: [`\u6399`].string() // U+6399 <cjk>
	0x58: utf32_to_str(0x22C24) // U+22C24 <cjk>
	0x59: [`\u6394`].string() // U+6394 <cjk>
	0x5A: [`\u63BD`].string() // U+63BD <cjk>
	0x5B: [`\u63F7`].string() // U+63F7 <cjk>
	0x5C: [`\u63D4`].string() // U+63D4 <cjk>
	0x5D: [`\u63D5`].string() // U+63D5 <cjk>
	0x5E: [`\u63DC`].string() // U+63DC <cjk>
	0x5F: [`\u63E0`].string() // U+63E0 <cjk>
	0x60: [`\u63EB`].string() // U+63EB <cjk>
	0x61: [`\u63EC`].string() // U+63EC <cjk>
	0x62: [`\u63F2`].string() // U+63F2 <cjk>
	0x63: [`\u6409`].string() // U+6409 <cjk>
	0x64: [`\u641E`].string() // U+641E <cjk>
	0x65: [`\u6425`].string() // U+6425 <cjk>
	0x66: [`\u6429`].string() // U+6429 <cjk>
	0x67: [`\u642F`].string() // U+642F <cjk>
	0x68: [`\u645A`].string() // U+645A <cjk>
	0x69: [`\u645B`].string() // U+645B <cjk>
	0x6A: [`\u645D`].string() // U+645D <cjk>
	0x6B: [`\u6473`].string() // U+6473 <cjk>
	0x6C: [`\u647D`].string() // U+647D <cjk>
	0x6D: [`\u6487`].string() // U+6487 <cjk>
	0x6E: [`\u6491`].string() // U+6491 <cjk>
	0x6F: [`\u649D`].string() // U+649D <cjk>
	0x70: [`\u649F`].string() // U+649F <cjk>
	0x71: [`\u64CB`].string() // U+64CB <cjk>
	0x72: [`\u64CC`].string() // U+64CC <cjk>
	0x73: [`\u64D5`].string() // U+64D5 <cjk>
	0x74: [`\u64D7`].string() // U+64D7 <cjk>
	0x75: utf32_to_str(0x22DE1) // U+22DE1 <cjk>
	0x76: [`\u64E4`].string() // U+64E4 <cjk>
	0x77: [`\u64E5`].string() // U+64E5 <cjk>
	0x78: [`\u64FF`].string() // U+64FF <cjk>
	0x79: [`\u6504`].string() // U+6504 <cjk>
	0x7A: [`\u3A6E`].string() // U+3A6E <cjk>
	0x7B: [`\u650F`].string() // U+650F <cjk>
	0x7C: [`\u6514`].string() // U+6514 <cjk>
	0x7D: [`\u6516`].string() // U+6516 <cjk>
	0x7E: [`\u3A73`].string() // U+3A73 <cjk>
	0x80: [`\u651E`].string() // U+651E <cjk>
	0x81: [`\u6532`].string() // U+6532 <cjk>
	0x82: [`\u6544`].string() // U+6544 <cjk>
	0x83: [`\u6554`].string() // U+6554 <cjk>
	0x84: [`\u656B`].string() // U+656B <cjk>
	0x85: [`\u657A`].string() // U+657A <cjk>
	0x86: [`\u6581`].string() // U+6581 <cjk>
	0x87: [`\u6584`].string() // U+6584 <cjk>
	0x88: [`\u6585`].string() // U+6585 <cjk>
	0x89: [`\u658A`].string() // U+658A <cjk>
	0x8A: [`\u65B2`].string() // U+65B2 <cjk>
	0x8B: [`\u65B5`].string() // U+65B5 <cjk>
	0x8C: [`\u65B8`].string() // U+65B8 <cjk>
	0x8D: [`\u65BF`].string() // U+65BF <cjk>
	0x8E: [`\u65C2`].string() // U+65C2 <cjk>
	0x8F: [`\u65C9`].string() // U+65C9 <cjk>
	0x90: [`\u65D4`].string() // U+65D4 <cjk>
	0x91: [`\u3AD6`].string() // U+3AD6 <cjk>
	0x92: [`\u65F2`].string() // U+65F2 <cjk>
	0x93: [`\u65F9`].string() // U+65F9 <cjk>
	0x94: [`\u65FC`].string() // U+65FC <cjk>
	0x95: [`\u6604`].string() // U+6604 <cjk>
	0x96: [`\u6608`].string() // U+6608 <cjk>
	0x97: [`\u6621`].string() // U+6621 <cjk>
	0x98: [`\u662A`].string() // U+662A <cjk>
	0x99: [`\u6645`].string() // U+6645 <cjk>
	0x9A: [`\u6651`].string() // U+6651 <cjk>
	0x9B: [`\u664E`].string() // U+664E <cjk>
	0x9C: [`\u3AEA`].string() // U+3AEA <cjk>
	0x9D: utf32_to_str(0x231C3) // U+231C3 <cjk>
	0x9E: [`\u6657`].string() // U+6657 <cjk>
	0x9F: [`\u665B`].string() // U+665B <cjk>
	0xA0: [`\u6663`].string() // U+6663 <cjk>
	0xA1: utf32_to_str(0x231F5) // U+231F5 <cjk>
	0xA2: utf32_to_str(0x231B6) // U+231B6 <cjk>
	0xA3: [`\u666A`].string() // U+666A <cjk>
	0xA4: [`\u666B`].string() // U+666B <cjk>
	0xA5: [`\u666C`].string() // U+666C <cjk>
	0xA6: [`\u666D`].string() // U+666D <cjk>
	0xA7: [`\u667B`].string() // U+667B <cjk>
	0xA8: [`\u6680`].string() // U+6680 <cjk>
	0xA9: [`\u6690`].string() // U+6690 <cjk>
	0xAA: [`\u6692`].string() // U+6692 <cjk>
	0xAB: [`\u6699`].string() // U+6699 <cjk>
	0xAC: [`\u3B0E`].string() // U+3B0E <cjk>
	0xAD: [`\u66AD`].string() // U+66AD <cjk>
	0xAE: [`\u66B1`].string() // U+66B1 <cjk>
	0xAF: [`\u66B5`].string() // U+66B5 <cjk>
	0xB0: [`\u3B1A`].string() // U+3B1A <cjk>
	0xB1: [`\u66BF`].string() // U+66BF <cjk>
	0xB2: [`\u3B1C`].string() // U+3B1C <cjk>
	0xB3: [`\u66EC`].string() // U+66EC <cjk>
	0xB4: [`\u3AD7`].string() // U+3AD7 <cjk>
	0xB5: [`\u6701`].string() // U+6701 <cjk>
	0xB6: [`\u6705`].string() // U+6705 <cjk>
	0xB7: [`\u6712`].string() // U+6712 <cjk>
	0xB8: utf32_to_str(0x23372) // U+23372 <cjk>
	0xB9: [`\u6719`].string() // U+6719 <cjk>
	0xBA: utf32_to_str(0x233D3) // U+233D3 <cjk>
	0xBB: utf32_to_str(0x233D2) // U+233D2 <cjk>
	0xBC: [`\u674C`].string() // U+674C <cjk>
	0xBD: [`\u674D`].string() // U+674D <cjk>
	0xBE: [`\u6754`].string() // U+6754 <cjk>
	0xBF: [`\u675D`].string() // U+675D <cjk>
	0xC0: utf32_to_str(0x233D0) // U+233D0 <cjk>
	0xC1: utf32_to_str(0x233E4) // U+233E4 <cjk>
	0xC2: utf32_to_str(0x233D5) // U+233D5 <cjk>
	0xC3: [`\u6774`].string() // U+6774 <cjk>
	0xC4: [`\u6776`].string() // U+6776 <cjk>
	0xC5: utf32_to_str(0x233DA) // U+233DA <cjk>
	0xC6: [`\u6792`].string() // U+6792 <cjk>
	0xC7: utf32_to_str(0x233DF) // U+233DF <cjk>
	0xC8: [`\u8363`].string() // U+8363 <cjk>
	0xC9: [`\u6810`].string() // U+6810 <cjk>
	0xCA: [`\u67B0`].string() // U+67B0 <cjk>
	0xCB: [`\u67B2`].string() // U+67B2 <cjk>
	0xCC: [`\u67C3`].string() // U+67C3 <cjk>
	0xCD: [`\u67C8`].string() // U+67C8 <cjk>
	0xCE: [`\u67D2`].string() // U+67D2 <cjk>
	0xCF: [`\u67D9`].string() // U+67D9 <cjk>
	0xD0: [`\u67DB`].string() // U+67DB <cjk>
	0xD1: [`\u67F0`].string() // U+67F0 <cjk>
	0xD2: [`\u67F7`].string() // U+67F7 <cjk>
	0xD3: utf32_to_str(0x2344A) // U+2344A <cjk>
	0xD4: utf32_to_str(0x23451) // U+23451 <cjk>
	0xD5: utf32_to_str(0x2344B) // U+2344B <cjk>
	0xD6: [`\u6818`].string() // U+6818 <cjk>
	0xD7: [`\u681F`].string() // U+681F <cjk>
	0xD8: [`\u682D`].string() // U+682D <cjk>
	0xD9: utf32_to_str(0x23465) // U+23465 <cjk>
	0xDA: [`\u6833`].string() // U+6833 <cjk>
	0xDB: [`\u683B`].string() // U+683B <cjk>
	0xDC: [`\u683E`].string() // U+683E <cjk>
	0xDD: [`\u6844`].string() // U+6844 <cjk>
	0xDE: [`\u6845`].string() // U+6845 <cjk>
	0xDF: [`\u6849`].string() // U+6849 <cjk>
	0xE0: [`\u684C`].string() // U+684C <cjk>
	0xE1: [`\u6855`].string() // U+6855 <cjk>
	0xE2: [`\u6857`].string() // U+6857 <cjk>
	0xE3: [`\u3B77`].string() // U+3B77 <cjk>
	0xE4: [`\u686B`].string() // U+686B <cjk>
	0xE5: [`\u686E`].string() // U+686E <cjk>
	0xE6: [`\u687A`].string() // U+687A <cjk>
	0xE7: [`\u687C`].string() // U+687C <cjk>
	0xE8: [`\u6882`].string() // U+6882 <cjk>
	0xE9: [`\u6890`].string() // U+6890 <cjk>
	0xEA: [`\u6896`].string() // U+6896 <cjk>
	0xEB: [`\u3B6D`].string() // U+3B6D <cjk>
	0xEC: [`\u6898`].string() // U+6898 <cjk>
	0xED: [`\u6899`].string() // U+6899 <cjk>
	0xEE: [`\u689A`].string() // U+689A <cjk>
	0xEF: [`\u689C`].string() // U+689C <cjk>
	0xF0: [`\u68AA`].string() // U+68AA <cjk>
	0xF1: [`\u68AB`].string() // U+68AB <cjk>
	0xF2: [`\u68B4`].string() // U+68B4 <cjk>
	0xF3: [`\u68BB`].string() // U+68BB <cjk>
	0xF4: [`\u68FB`].string() // U+68FB <cjk>
	0xF5: utf32_to_str(0x234E4) // U+234E4 <cjk>
	0xF6: utf32_to_str(0x2355A) // U+2355A <cjk>
	0xF7: [`\uFA13`].string() // U+FA13 CJK COMPATIBILITY IDEOGRAPH-FA13
	0xF8: [`\u68C3`].string() // U+68C3 <cjk>
	0xF9: [`\u68C5`].string() // U+68C5 <cjk>
	0xFA: [`\u68CC`].string() // U+68CC <cjk>
	0xFB: [`\u68CF`].string() // U+68CF <cjk>
	0xFC: [`\u68D6`].string() // U+68D6 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xe2 = {
	0x40: [`\u78E7`].string() // U+78E7 <cjk>
	0x41: [`\u78DA`].string() // U+78DA <cjk>
	0x42: [`\u78FD`].string() // U+78FD <cjk>
	0x43: [`\u78F4`].string() // U+78F4 <cjk>
	0x44: [`\u7907`].string() // U+7907 <cjk>
	0x45: [`\u7912`].string() // U+7912 <cjk>
	0x46: [`\u7911`].string() // U+7911 <cjk>
	0x47: [`\u7919`].string() // U+7919 <cjk>
	0x48: [`\u792C`].string() // U+792C <cjk>
	0x49: [`\u792B`].string() // U+792B <cjk>
	0x4A: [`\u7940`].string() // U+7940 <cjk>
	0x4B: [`\u7960`].string() // U+7960 <cjk>
	0x4C: [`\u7957`].string() // U+7957 <cjk>
	0x4D: [`\u795F`].string() // U+795F <cjk>
	0x4E: [`\u795A`].string() // U+795A <cjk>
	0x4F: [`\u7955`].string() // U+7955 <cjk>
	0x50: [`\u7953`].string() // U+7953 <cjk>
	0x51: [`\u797A`].string() // U+797A <cjk>
	0x52: [`\u797F`].string() // U+797F <cjk>
	0x53: [`\u798A`].string() // U+798A <cjk>
	0x54: [`\u799D`].string() // U+799D <cjk>
	0x55: [`\u79A7`].string() // U+79A7 <cjk>
	0x56: [`\u9F4B`].string() // U+9F4B <cjk>
	0x57: [`\u79AA`].string() // U+79AA <cjk>
	0x58: [`\u79AE`].string() // U+79AE <cjk>
	0x59: [`\u79B3`].string() // U+79B3 <cjk>
	0x5A: [`\u79B9`].string() // U+79B9 <cjk>
	0x5B: [`\u79BA`].string() // U+79BA <cjk>
	0x5C: [`\u79C9`].string() // U+79C9 <cjk>
	0x5D: [`\u79D5`].string() // U+79D5 <cjk>
	0x5E: [`\u79E7`].string() // U+79E7 <cjk>
	0x5F: [`\u79EC`].string() // U+79EC <cjk>
	0x60: [`\u79E1`].string() // U+79E1 <cjk>
	0x61: [`\u79E3`].string() // U+79E3 <cjk>
	0x62: [`\u7A08`].string() // U+7A08 <cjk>
	0x63: [`\u7A0D`].string() // U+7A0D <cjk>
	0x64: [`\u7A18`].string() // U+7A18 <cjk>
	0x65: [`\u7A19`].string() // U+7A19 <cjk>
	0x66: [`\u7A20`].string() // U+7A20 <cjk>
	0x67: [`\u7A1F`].string() // U+7A1F <cjk>
	0x68: [`\u7980`].string() // U+7980 <cjk>
	0x69: [`\u7A31`].string() // U+7A31 <cjk>
	0x6A: [`\u7A3B`].string() // U+7A3B <cjk>
	0x6B: [`\u7A3E`].string() // U+7A3E <cjk>
	0x6C: [`\u7A37`].string() // U+7A37 <cjk>
	0x6D: [`\u7A43`].string() // U+7A43 <cjk>
	0x6E: [`\u7A57`].string() // U+7A57 <cjk>
	0x6F: [`\u7A49`].string() // U+7A49 <cjk>
	0x70: [`\u7A61`].string() // U+7A61 <cjk>
	0x71: [`\u7A62`].string() // U+7A62 <cjk>
	0x72: [`\u7A69`].string() // U+7A69 <cjk>
	0x73: [`\u9F9D`].string() // U+9F9D <cjk>
	0x74: [`\u7A70`].string() // U+7A70 <cjk>
	0x75: [`\u7A79`].string() // U+7A79 <cjk>
	0x76: [`\u7A7D`].string() // U+7A7D <cjk>
	0x77: [`\u7A88`].string() // U+7A88 <cjk>
	0x78: [`\u7A97`].string() // U+7A97 <cjk>
	0x79: [`\u7A95`].string() // U+7A95 <cjk>
	0x7A: [`\u7A98`].string() // U+7A98 <cjk>
	0x7B: [`\u7A96`].string() // U+7A96 <cjk>
	0x7C: [`\u7AA9`].string() // U+7AA9 <cjk>
	0x7D: [`\u7AC8`].string() // U+7AC8 <cjk>
	0x7E: [`\u7AB0`].string() // U+7AB0 <cjk>
	0x80: [`\u7AB6`].string() // U+7AB6 <cjk>
	0x81: [`\u7AC5`].string() // U+7AC5 <cjk>
	0x82: [`\u7AC4`].string() // U+7AC4 <cjk>
	0x83: [`\u7ABF`].string() // U+7ABF <cjk>
	0x84: [`\u9083`].string() // U+9083 <cjk>
	0x85: [`\u7AC7`].string() // U+7AC7 <cjk>
	0x86: [`\u7ACA`].string() // U+7ACA <cjk>
	0x87: [`\u7ACD`].string() // U+7ACD <cjk>
	0x88: [`\u7ACF`].string() // U+7ACF <cjk>
	0x89: [`\u7AD5`].string() // U+7AD5 <cjk>
	0x8A: [`\u7AD3`].string() // U+7AD3 <cjk>
	0x8B: [`\u7AD9`].string() // U+7AD9 <cjk>
	0x8C: [`\u7ADA`].string() // U+7ADA <cjk>
	0x8D: [`\u7ADD`].string() // U+7ADD <cjk>
	0x8E: [`\u7AE1`].string() // U+7AE1 <cjk>
	0x8F: [`\u7AE2`].string() // U+7AE2 <cjk>
	0x90: [`\u7AE6`].string() // U+7AE6 <cjk>
	0x91: [`\u7AED`].string() // U+7AED <cjk>
	0x92: [`\u7AF0`].string() // U+7AF0 <cjk>
	0x93: [`\u7B02`].string() // U+7B02 <cjk>
	0x94: [`\u7B0F`].string() // U+7B0F <cjk>
	0x95: [`\u7B0A`].string() // U+7B0A <cjk>
	0x96: [`\u7B06`].string() // U+7B06 <cjk>
	0x97: [`\u7B33`].string() // U+7B33 <cjk>
	0x98: [`\u7B18`].string() // U+7B18 <cjk>
	0x99: [`\u7B19`].string() // U+7B19 <cjk>
	0x9A: [`\u7B1E`].string() // U+7B1E <cjk>
	0x9B: [`\u7B35`].string() // U+7B35 <cjk>
	0x9C: [`\u7B28`].string() // U+7B28 <cjk>
	0x9D: [`\u7B36`].string() // U+7B36 <cjk>
	0x9E: [`\u7B50`].string() // U+7B50 <cjk>
	0x9F: [`\u7B7A`].string() // U+7B7A <cjk>
	0xA0: [`\u7B04`].string() // U+7B04 <cjk>
	0xA1: [`\u7B4D`].string() // U+7B4D <cjk>
	0xA2: [`\u7B0B`].string() // U+7B0B <cjk>
	0xA3: [`\u7B4C`].string() // U+7B4C <cjk>
	0xA4: [`\u7B45`].string() // U+7B45 <cjk>
	0xA5: [`\u7B75`].string() // U+7B75 <cjk>
	0xA6: [`\u7B65`].string() // U+7B65 <cjk>
	0xA7: [`\u7B74`].string() // U+7B74 <cjk>
	0xA8: [`\u7B67`].string() // U+7B67 <cjk>
	0xA9: [`\u7B70`].string() // U+7B70 <cjk>
	0xAA: [`\u7B71`].string() // U+7B71 <cjk>
	0xAB: [`\u7B6C`].string() // U+7B6C <cjk>
	0xAC: [`\u7B6E`].string() // U+7B6E <cjk>
	0xAD: [`\u7B9D`].string() // U+7B9D <cjk>
	0xAE: [`\u7B98`].string() // U+7B98 <cjk>
	0xAF: [`\u7B9F`].string() // U+7B9F <cjk>
	0xB0: [`\u7B8D`].string() // U+7B8D <cjk>
	0xB1: [`\u7B9C`].string() // U+7B9C <cjk>
	0xB2: [`\u7B9A`].string() // U+7B9A <cjk>
	0xB3: [`\u7B8B`].string() // U+7B8B <cjk>
	0xB4: [`\u7B92`].string() // U+7B92 <cjk>
	0xB5: [`\u7B8F`].string() // U+7B8F <cjk>
	0xB6: [`\u7B5D`].string() // U+7B5D <cjk>
	0xB7: [`\u7B99`].string() // U+7B99 <cjk>
	0xB8: [`\u7BCB`].string() // U+7BCB <cjk>
	0xB9: [`\u7BC1`].string() // U+7BC1 <cjk>
	0xBA: [`\u7BCC`].string() // U+7BCC <cjk>
	0xBB: [`\u7BCF`].string() // U+7BCF <cjk>
	0xBC: [`\u7BB4`].string() // U+7BB4 <cjk>
	0xBD: [`\u7BC6`].string() // U+7BC6 <cjk>
	0xBE: [`\u7BDD`].string() // U+7BDD <cjk>
	0xBF: [`\u7BE9`].string() // U+7BE9 <cjk>
	0xC0: [`\u7C11`].string() // U+7C11 <cjk>
	0xC1: [`\u7C14`].string() // U+7C14 <cjk>
	0xC2: [`\u7BE6`].string() // U+7BE6 <cjk>
	0xC3: [`\u7BE5`].string() // U+7BE5 <cjk>
	0xC4: [`\u7C60`].string() // U+7C60 <cjk>
	0xC5: [`\u7C00`].string() // U+7C00 <cjk>
	0xC6: [`\u7C07`].string() // U+7C07 <cjk>
	0xC7: [`\u7C13`].string() // U+7C13 <cjk>
	0xC8: [`\u7BF3`].string() // U+7BF3 <cjk>
	0xC9: [`\u7BF7`].string() // U+7BF7 <cjk>
	0xCA: [`\u7C17`].string() // U+7C17 <cjk>
	0xCB: [`\u7C0D`].string() // U+7C0D <cjk>
	0xCC: [`\u7BF6`].string() // U+7BF6 <cjk>
	0xCD: [`\u7C23`].string() // U+7C23 <cjk>
	0xCE: [`\u7C27`].string() // U+7C27 <cjk>
	0xCF: [`\u7C2A`].string() // U+7C2A <cjk>
	0xD0: [`\u7C1F`].string() // U+7C1F <cjk>
	0xD1: [`\u7C37`].string() // U+7C37 <cjk>
	0xD2: [`\u7C2B`].string() // U+7C2B <cjk>
	0xD3: [`\u7C3D`].string() // U+7C3D <cjk>
	0xD4: [`\u7C4C`].string() // U+7C4C <cjk>
	0xD5: [`\u7C43`].string() // U+7C43 <cjk>
	0xD6: [`\u7C54`].string() // U+7C54 <cjk>
	0xD7: [`\u7C4F`].string() // U+7C4F <cjk>
	0xD8: [`\u7C40`].string() // U+7C40 <cjk>
	0xD9: [`\u7C50`].string() // U+7C50 <cjk>
	0xDA: [`\u7C58`].string() // U+7C58 <cjk>
	0xDB: [`\u7C5F`].string() // U+7C5F <cjk>
	0xDC: [`\u7C64`].string() // U+7C64 <cjk>
	0xDD: [`\u7C56`].string() // U+7C56 <cjk>
	0xDE: [`\u7C65`].string() // U+7C65 <cjk>
	0xDF: [`\u7C6C`].string() // U+7C6C <cjk>
	0xE0: [`\u7C75`].string() // U+7C75 <cjk>
	0xE1: [`\u7C83`].string() // U+7C83 <cjk>
	0xE2: [`\u7C90`].string() // U+7C90 <cjk>
	0xE3: [`\u7CA4`].string() // U+7CA4 <cjk>
	0xE4: [`\u7CAD`].string() // U+7CAD <cjk>
	0xE5: [`\u7CA2`].string() // U+7CA2 <cjk>
	0xE6: [`\u7CAB`].string() // U+7CAB <cjk>
	0xE7: [`\u7CA1`].string() // U+7CA1 <cjk>
	0xE8: [`\u7CA8`].string() // U+7CA8 <cjk>
	0xE9: [`\u7CB3`].string() // U+7CB3 <cjk>
	0xEA: [`\u7CB2`].string() // U+7CB2 <cjk>
	0xEB: [`\u7CB1`].string() // U+7CB1 <cjk>
	0xEC: [`\u7CAE`].string() // U+7CAE <cjk>
	0xED: [`\u7CB9`].string() // U+7CB9 <cjk>
	0xEE: [`\u7CBD`].string() // U+7CBD <cjk>
	0xEF: [`\u7CC0`].string() // U+7CC0 <cjk>
	0xF0: [`\u7CC5`].string() // U+7CC5 <cjk>
	0xF1: [`\u7CC2`].string() // U+7CC2 <cjk>
	0xF2: [`\u7CD8`].string() // U+7CD8 <cjk>
	0xF3: [`\u7CD2`].string() // U+7CD2 <cjk>
	0xF4: [`\u7CDC`].string() // U+7CDC <cjk>
	0xF5: [`\u7CE2`].string() // U+7CE2 <cjk>
	0xF6: [`\u9B3B`].string() // U+9B3B <cjk>
	0xF7: [`\u7CEF`].string() // U+7CEF <cjk>
	0xF8: [`\u7CF2`].string() // U+7CF2 <cjk>
	0xF9: [`\u7CF4`].string() // U+7CF4 <cjk>
	0xFA: [`\u7CF6`].string() // U+7CF6 <cjk>
	0xFB: [`\u7CFA`].string() // U+7CFA <cjk>
	0xFC: [`\u7D06`].string() // U+7D06 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x9a = {
	0x40: [`\u54AB`].string() // U+54AB <cjk>
	0x41: [`\u54C2`].string() // U+54C2 <cjk>
	0x42: [`\u54A4`].string() // U+54A4 <cjk>
	0x43: [`\u54BE`].string() // U+54BE <cjk>
	0x44: [`\u54BC`].string() // U+54BC <cjk>
	0x45: [`\u54D8`].string() // U+54D8 <cjk>
	0x46: [`\u54E5`].string() // U+54E5 <cjk>
	0x47: [`\u54E6`].string() // U+54E6 <cjk>
	0x48: [`\u550F`].string() // U+550F <cjk>
	0x49: [`\u5514`].string() // U+5514 <cjk>
	0x4A: [`\u54FD`].string() // U+54FD <cjk>
	0x4B: [`\u54EE`].string() // U+54EE <cjk>
	0x4C: [`\u54ED`].string() // U+54ED <cjk>
	0x4D: [`\u54FA`].string() // U+54FA <cjk>
	0x4E: [`\u54E2`].string() // U+54E2 <cjk>
	0x4F: [`\u5539`].string() // U+5539 <cjk>
	0x50: [`\u5540`].string() // U+5540 <cjk>
	0x51: [`\u5563`].string() // U+5563 <cjk>
	0x52: [`\u554C`].string() // U+554C <cjk>
	0x53: [`\u552E`].string() // U+552E <cjk>
	0x54: [`\u555C`].string() // U+555C <cjk>
	0x55: [`\u5545`].string() // U+5545 <cjk>
	0x56: [`\u5556`].string() // U+5556 <cjk>
	0x57: [`\u5557`].string() // U+5557 <cjk>
	0x58: [`\u5538`].string() // U+5538 <cjk>
	0x59: [`\u5533`].string() // U+5533 <cjk>
	0x5A: [`\u555D`].string() // U+555D <cjk>
	0x5B: [`\u5599`].string() // U+5599 <cjk>
	0x5C: [`\u5580`].string() // U+5580 <cjk>
	0x5D: [`\u54AF`].string() // U+54AF <cjk>
	0x5E: [`\u558A`].string() // U+558A <cjk>
	0x5F: [`\u559F`].string() // U+559F <cjk>
	0x60: [`\u557B`].string() // U+557B <cjk>
	0x61: [`\u557E`].string() // U+557E <cjk>
	0x62: [`\u5598`].string() // U+5598 <cjk>
	0x63: [`\u559E`].string() // U+559E <cjk>
	0x64: [`\u55AE`].string() // U+55AE <cjk>
	0x65: [`\u557C`].string() // U+557C <cjk>
	0x66: [`\u5583`].string() // U+5583 <cjk>
	0x67: [`\u55A9`].string() // U+55A9 <cjk>
	0x68: [`\u5587`].string() // U+5587 <cjk>
	0x69: [`\u55A8`].string() // U+55A8 <cjk>
	0x6A: [`\u55DA`].string() // U+55DA <cjk>
	0x6B: [`\u55C5`].string() // U+55C5 <cjk>
	0x6C: [`\u55DF`].string() // U+55DF <cjk>
	0x6D: [`\u55C4`].string() // U+55C4 <cjk>
	0x6E: [`\u55DC`].string() // U+55DC <cjk>
	0x6F: [`\u55E4`].string() // U+55E4 <cjk>
	0x70: [`\u55D4`].string() // U+55D4 <cjk>
	0x71: [`\u5614`].string() // U+5614 <cjk>
	0x72: [`\u55F7`].string() // U+55F7 <cjk>
	0x73: [`\u5616`].string() // U+5616 <cjk>
	0x74: [`\u55FE`].string() // U+55FE <cjk>
	0x75: [`\u55FD`].string() // U+55FD <cjk>
	0x76: [`\u561B`].string() // U+561B <cjk>
	0x77: [`\u55F9`].string() // U+55F9 <cjk>
	0x78: [`\u564E`].string() // U+564E <cjk>
	0x79: [`\u5650`].string() // U+5650 <cjk>
	0x7A: [`\u71DF`].string() // U+71DF <cjk>
	0x7B: [`\u5634`].string() // U+5634 <cjk>
	0x7C: [`\u5636`].string() // U+5636 <cjk>
	0x7D: [`\u5632`].string() // U+5632 <cjk>
	0x7E: [`\u5638`].string() // U+5638 <cjk>
	0x80: [`\u566B`].string() // U+566B <cjk>
	0x81: [`\u5664`].string() // U+5664 <cjk>
	0x82: [`\u562F`].string() // U+562F <cjk>
	0x83: [`\u566C`].string() // U+566C <cjk>
	0x84: [`\u566A`].string() // U+566A <cjk>
	0x85: [`\u5686`].string() // U+5686 <cjk>
	0x86: [`\u5680`].string() // U+5680 <cjk>
	0x87: [`\u568A`].string() // U+568A <cjk>
	0x88: [`\u56A0`].string() // U+56A0 <cjk>
	0x89: [`\u5694`].string() // U+5694 <cjk>
	0x8A: [`\u568F`].string() // U+568F <cjk>
	0x8B: [`\u56A5`].string() // U+56A5 <cjk>
	0x8C: [`\u56AE`].string() // U+56AE <cjk>
	0x8D: [`\u56B6`].string() // U+56B6 <cjk>
	0x8E: [`\u56B4`].string() // U+56B4 <cjk>
	0x8F: [`\u56C2`].string() // U+56C2 <cjk>
	0x90: [`\u56BC`].string() // U+56BC <cjk>
	0x91: [`\u56C1`].string() // U+56C1 <cjk>
	0x92: [`\u56C3`].string() // U+56C3 <cjk>
	0x93: [`\u56C0`].string() // U+56C0 <cjk>
	0x94: [`\u56C8`].string() // U+56C8 <cjk>
	0x95: [`\u56CE`].string() // U+56CE <cjk>
	0x96: [`\u56D1`].string() // U+56D1 <cjk>
	0x97: [`\u56D3`].string() // U+56D3 <cjk>
	0x98: [`\u56D7`].string() // U+56D7 <cjk>
	0x99: [`\u56EE`].string() // U+56EE <cjk>
	0x9A: [`\u56F9`].string() // U+56F9 <cjk>
	0x9B: [`\u5700`].string() // U+5700 <cjk>
	0x9C: [`\u56FF`].string() // U+56FF <cjk>
	0x9D: [`\u5704`].string() // U+5704 <cjk>
	0x9E: [`\u5709`].string() // U+5709 <cjk>
	0x9F: [`\u5708`].string() // U+5708 <cjk>
	0xA0: [`\u570B`].string() // U+570B <cjk>
	0xA1: [`\u570D`].string() // U+570D <cjk>
	0xA2: [`\u5713`].string() // U+5713 <cjk>
	0xA3: [`\u5718`].string() // U+5718 <cjk>
	0xA4: [`\u5716`].string() // U+5716 <cjk>
	0xA5: [`\u55C7`].string() // U+55C7 <cjk>
	0xA6: [`\u571C`].string() // U+571C <cjk>
	0xA7: [`\u5726`].string() // U+5726 <cjk>
	0xA8: [`\u5737`].string() // U+5737 <cjk>
	0xA9: [`\u5738`].string() // U+5738 <cjk>
	0xAA: [`\u574E`].string() // U+574E <cjk>
	0xAB: [`\u573B`].string() // U+573B <cjk>
	0xAC: [`\u5740`].string() // U+5740 <cjk>
	0xAD: [`\u574F`].string() // U+574F <cjk>
	0xAE: [`\u5769`].string() // U+5769 <cjk>
	0xAF: [`\u57C0`].string() // U+57C0 <cjk>
	0xB0: [`\u5788`].string() // U+5788 <cjk>
	0xB1: [`\u5761`].string() // U+5761 <cjk>
	0xB2: [`\u577F`].string() // U+577F <cjk>
	0xB3: [`\u5789`].string() // U+5789 <cjk>
	0xB4: [`\u5793`].string() // U+5793 <cjk>
	0xB5: [`\u57A0`].string() // U+57A0 <cjk>
	0xB6: [`\u57B3`].string() // U+57B3 <cjk>
	0xB7: [`\u57A4`].string() // U+57A4 <cjk>
	0xB8: [`\u57AA`].string() // U+57AA <cjk>
	0xB9: [`\u57B0`].string() // U+57B0 <cjk>
	0xBA: [`\u57C3`].string() // U+57C3 <cjk>
	0xBB: [`\u57C6`].string() // U+57C6 <cjk>
	0xBC: [`\u57D4`].string() // U+57D4 <cjk>
	0xBD: [`\u57D2`].string() // U+57D2 <cjk>
	0xBE: [`\u57D3`].string() // U+57D3 <cjk>
	0xBF: [`\u580A`].string() // U+580A <cjk>
	0xC0: [`\u57D6`].string() // U+57D6 <cjk>
	0xC1: [`\u57E3`].string() // U+57E3 <cjk>
	0xC2: [`\u580B`].string() // U+580B <cjk>
	0xC3: [`\u5819`].string() // U+5819 <cjk>
	0xC4: [`\u581D`].string() // U+581D <cjk>
	0xC5: [`\u5872`].string() // U+5872 <cjk>
	0xC6: [`\u5821`].string() // U+5821 <cjk>
	0xC7: [`\u5862`].string() // U+5862 <cjk>
	0xC8: [`\u584B`].string() // U+584B <cjk>
	0xC9: [`\u5870`].string() // U+5870 <cjk>
	0xCA: [`\u6BC0`].string() // U+6BC0 <cjk>
	0xCB: [`\u5852`].string() // U+5852 <cjk>
	0xCC: [`\u583D`].string() // U+583D <cjk>
	0xCD: [`\u5879`].string() // U+5879 <cjk>
	0xCE: [`\u5885`].string() // U+5885 <cjk>
	0xCF: [`\u58B9`].string() // U+58B9 <cjk>
	0xD0: [`\u589F`].string() // U+589F <cjk>
	0xD1: [`\u58AB`].string() // U+58AB <cjk>
	0xD2: [`\u58BA`].string() // U+58BA <cjk>
	0xD3: [`\u58DE`].string() // U+58DE <cjk>
	0xD4: [`\u58BB`].string() // U+58BB <cjk>
	0xD5: [`\u58B8`].string() // U+58B8 <cjk>
	0xD6: [`\u58AE`].string() // U+58AE <cjk>
	0xD7: [`\u58C5`].string() // U+58C5 <cjk>
	0xD8: [`\u58D3`].string() // U+58D3 <cjk>
	0xD9: [`\u58D1`].string() // U+58D1 <cjk>
	0xDA: [`\u58D7`].string() // U+58D7 <cjk>
	0xDB: [`\u58D9`].string() // U+58D9 <cjk>
	0xDC: [`\u58D8`].string() // U+58D8 <cjk>
	0xDD: [`\u58E5`].string() // U+58E5 <cjk>
	0xDE: [`\u58DC`].string() // U+58DC <cjk>
	0xDF: [`\u58E4`].string() // U+58E4 <cjk>
	0xE0: [`\u58DF`].string() // U+58DF <cjk>
	0xE1: [`\u58EF`].string() // U+58EF <cjk>
	0xE2: [`\u58FA`].string() // U+58FA <cjk>
	0xE3: [`\u58F9`].string() // U+58F9 <cjk>
	0xE4: [`\u58FB`].string() // U+58FB <cjk>
	0xE5: [`\u58FC`].string() // U+58FC <cjk>
	0xE6: [`\u58FD`].string() // U+58FD <cjk>
	0xE7: [`\u5902`].string() // U+5902 <cjk>
	0xE8: [`\u590A`].string() // U+590A <cjk>
	0xE9: [`\u5910`].string() // U+5910 <cjk>
	0xEA: [`\u591B`].string() // U+591B <cjk>
	0xEB: [`\u68A6`].string() // U+68A6 <cjk>
	0xEC: [`\u5925`].string() // U+5925 <cjk>
	0xED: [`\u592C`].string() // U+592C <cjk>
	0xEE: [`\u592D`].string() // U+592D <cjk>
	0xEF: [`\u5932`].string() // U+5932 <cjk>
	0xF0: [`\u5938`].string() // U+5938 <cjk>
	0xF1: [`\u593E`].string() // U+593E <cjk>
	0xF2: [`\u7AD2`].string() // U+7AD2 <cjk>
	0xF3: [`\u5955`].string() // U+5955 <cjk>
	0xF4: [`\u5950`].string() // U+5950 <cjk>
	0xF5: [`\u594E`].string() // U+594E <cjk>
	0xF6: [`\u595A`].string() // U+595A <cjk>
	0xF7: [`\u5958`].string() // U+5958 <cjk>
	0xF8: [`\u5962`].string() // U+5962 <cjk>
	0xF9: [`\u5960`].string() // U+5960 <cjk>
	0xFA: [`\u5967`].string() // U+5967 <cjk>
	0xFB: [`\u596C`].string() // U+596C <cjk>
	0xFC: [`\u5969`].string() // U+5969 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xe5 = {
	0x40: [`\u8541`].string() // U+8541 <cjk>
	0x41: [`\u8602`].string() // U+8602 <cjk>
	0x42: [`\u854B`].string() // U+854B <cjk>
	0x43: [`\u8555`].string() // U+8555 <cjk>
	0x44: [`\u8580`].string() // U+8580 <cjk>
	0x45: [`\u85A4`].string() // U+85A4 <cjk>
	0x46: [`\u8588`].string() // U+8588 <cjk>
	0x47: [`\u8591`].string() // U+8591 <cjk>
	0x48: [`\u858A`].string() // U+858A <cjk>
	0x49: [`\u85A8`].string() // U+85A8 <cjk>
	0x4A: [`\u856D`].string() // U+856D <cjk>
	0x4B: [`\u8594`].string() // U+8594 <cjk>
	0x4C: [`\u859B`].string() // U+859B <cjk>
	0x4D: [`\u85EA`].string() // U+85EA <cjk>
	0x4E: [`\u8587`].string() // U+8587 <cjk>
	0x4F: [`\u859C`].string() // U+859C <cjk>
	0x50: [`\u8577`].string() // U+8577 <cjk>
	0x51: [`\u857E`].string() // U+857E <cjk>
	0x52: [`\u8590`].string() // U+8590 <cjk>
	0x53: [`\u85C9`].string() // U+85C9 <cjk>
	0x54: [`\u85BA`].string() // U+85BA <cjk>
	0x55: [`\u85CF`].string() // U+85CF <cjk>
	0x56: [`\u85B9`].string() // U+85B9 <cjk>
	0x57: [`\u85D0`].string() // U+85D0 <cjk>
	0x58: [`\u85D5`].string() // U+85D5 <cjk>
	0x59: [`\u85DD`].string() // U+85DD <cjk>
	0x5A: [`\u85E5`].string() // U+85E5 <cjk>
	0x5B: [`\u85DC`].string() // U+85DC <cjk>
	0x5C: [`\u85F9`].string() // U+85F9 <cjk>
	0x5D: [`\u860A`].string() // U+860A <cjk>
	0x5E: [`\u8613`].string() // U+8613 <cjk>
	0x5F: [`\u860B`].string() // U+860B <cjk>
	0x60: [`\u85FE`].string() // U+85FE <cjk>
	0x61: [`\u85FA`].string() // U+85FA <cjk>
	0x62: [`\u8606`].string() // U+8606 <cjk>
	0x63: [`\u8622`].string() // U+8622 <cjk>
	0x64: [`\u861A`].string() // U+861A <cjk>
	0x65: [`\u8630`].string() // U+8630 <cjk>
	0x66: [`\u863F`].string() // U+863F <cjk>
	0x67: [`\u864D`].string() // U+864D <cjk>
	0x68: [`\u4E55`].string() // U+4E55 <cjk>
	0x69: [`\u8654`].string() // U+8654 <cjk>
	0x6A: [`\u865F`].string() // U+865F <cjk>
	0x6B: [`\u8667`].string() // U+8667 <cjk>
	0x6C: [`\u8671`].string() // U+8671 <cjk>
	0x6D: [`\u8693`].string() // U+8693 <cjk>
	0x6E: [`\u86A3`].string() // U+86A3 <cjk>
	0x6F: [`\u86A9`].string() // U+86A9 <cjk>
	0x70: [`\u86AA`].string() // U+86AA <cjk>
	0x71: [`\u868B`].string() // U+868B <cjk>
	0x72: [`\u868C`].string() // U+868C <cjk>
	0x73: [`\u86B6`].string() // U+86B6 <cjk>
	0x74: [`\u86AF`].string() // U+86AF <cjk>
	0x75: [`\u86C4`].string() // U+86C4 <cjk>
	0x76: [`\u86C6`].string() // U+86C6 <cjk>
	0x77: [`\u86B0`].string() // U+86B0 <cjk>
	0x78: [`\u86C9`].string() // U+86C9 <cjk>
	0x79: [`\u8823`].string() // U+8823 <cjk>
	0x7A: [`\u86AB`].string() // U+86AB <cjk>
	0x7B: [`\u86D4`].string() // U+86D4 <cjk>
	0x7C: [`\u86DE`].string() // U+86DE <cjk>
	0x7D: [`\u86E9`].string() // U+86E9 <cjk>
	0x7E: [`\u86EC`].string() // U+86EC <cjk>
	0x80: [`\u86DF`].string() // U+86DF <cjk>
	0x81: [`\u86DB`].string() // U+86DB <cjk>
	0x82: [`\u86EF`].string() // U+86EF <cjk>
	0x83: [`\u8712`].string() // U+8712 <cjk>
	0x84: [`\u8706`].string() // U+8706 <cjk>
	0x85: [`\u8708`].string() // U+8708 <cjk>
	0x86: [`\u8700`].string() // U+8700 <cjk>
	0x87: [`\u8703`].string() // U+8703 <cjk>
	0x88: [`\u86FB`].string() // U+86FB <cjk>
	0x89: [`\u8711`].string() // U+8711 <cjk>
	0x8A: [`\u8709`].string() // U+8709 <cjk>
	0x8B: [`\u870D`].string() // U+870D <cjk>
	0x8C: [`\u86F9`].string() // U+86F9 <cjk>
	0x8D: [`\u870A`].string() // U+870A <cjk>
	0x8E: [`\u8734`].string() // U+8734 <cjk>
	0x8F: [`\u873F`].string() // U+873F <cjk>
	0x90: [`\u8737`].string() // U+8737 <cjk>
	0x91: [`\u873B`].string() // U+873B <cjk>
	0x92: [`\u8725`].string() // U+8725 <cjk>
	0x93: [`\u8729`].string() // U+8729 <cjk>
	0x94: [`\u871A`].string() // U+871A <cjk>
	0x95: [`\u8760`].string() // U+8760 <cjk>
	0x96: [`\u875F`].string() // U+875F <cjk>
	0x97: [`\u8778`].string() // U+8778 <cjk>
	0x98: [`\u874C`].string() // U+874C <cjk>
	0x99: [`\u874E`].string() // U+874E <cjk>
	0x9A: [`\u8774`].string() // U+8774 <cjk>
	0x9B: [`\u8757`].string() // U+8757 <cjk>
	0x9C: [`\u8768`].string() // U+8768 <cjk>
	0x9D: [`\u876E`].string() // U+876E <cjk>
	0x9E: [`\u8759`].string() // U+8759 <cjk>
	0x9F: [`\u8753`].string() // U+8753 <cjk>
	0xA0: [`\u8763`].string() // U+8763 <cjk>
	0xA1: [`\u876A`].string() // U+876A <cjk>
	0xA2: [`\u8805`].string() // U+8805 <cjk>
	0xA3: [`\u87A2`].string() // U+87A2 <cjk>
	0xA4: [`\u879F`].string() // U+879F <cjk>
	0xA5: [`\u8782`].string() // U+8782 <cjk>
	0xA6: [`\u87AF`].string() // U+87AF <cjk>
	0xA7: [`\u87CB`].string() // U+87CB <cjk>
	0xA8: [`\u87BD`].string() // U+87BD <cjk>
	0xA9: [`\u87C0`].string() // U+87C0 <cjk>
	0xAA: [`\u87D0`].string() // U+87D0 <cjk>
	0xAB: [`\u96D6`].string() // U+96D6 <cjk>
	0xAC: [`\u87AB`].string() // U+87AB <cjk>
	0xAD: [`\u87C4`].string() // U+87C4 <cjk>
	0xAE: [`\u87B3`].string() // U+87B3 <cjk>
	0xAF: [`\u87C7`].string() // U+87C7 <cjk>
	0xB0: [`\u87C6`].string() // U+87C6 <cjk>
	0xB1: [`\u87BB`].string() // U+87BB <cjk>
	0xB2: [`\u87EF`].string() // U+87EF <cjk>
	0xB3: [`\u87F2`].string() // U+87F2 <cjk>
	0xB4: [`\u87E0`].string() // U+87E0 <cjk>
	0xB5: [`\u880F`].string() // U+880F <cjk>
	0xB6: [`\u880D`].string() // U+880D <cjk>
	0xB7: [`\u87FE`].string() // U+87FE <cjk>
	0xB8: [`\u87F6`].string() // U+87F6 <cjk>
	0xB9: [`\u87F7`].string() // U+87F7 <cjk>
	0xBA: [`\u880E`].string() // U+880E <cjk>
	0xBB: [`\u87D2`].string() // U+87D2 <cjk>
	0xBC: [`\u8811`].string() // U+8811 <cjk>
	0xBD: [`\u8816`].string() // U+8816 <cjk>
	0xBE: [`\u8815`].string() // U+8815 <cjk>
	0xBF: [`\u8822`].string() // U+8822 <cjk>
	0xC0: [`\u8821`].string() // U+8821 <cjk>
	0xC1: [`\u8831`].string() // U+8831 <cjk>
	0xC2: [`\u8836`].string() // U+8836 <cjk>
	0xC3: [`\u8839`].string() // U+8839 <cjk>
	0xC4: [`\u8827`].string() // U+8827 <cjk>
	0xC5: [`\u883B`].string() // U+883B <cjk>
	0xC6: [`\u8844`].string() // U+8844 <cjk>
	0xC7: [`\u8842`].string() // U+8842 <cjk>
	0xC8: [`\u8852`].string() // U+8852 <cjk>
	0xC9: [`\u8859`].string() // U+8859 <cjk>
	0xCA: [`\u885E`].string() // U+885E <cjk>
	0xCB: [`\u8862`].string() // U+8862 <cjk>
	0xCC: [`\u886B`].string() // U+886B <cjk>
	0xCD: [`\u8881`].string() // U+8881 <cjk>
	0xCE: [`\u887E`].string() // U+887E <cjk>
	0xCF: [`\u889E`].string() // U+889E <cjk>
	0xD0: [`\u8875`].string() // U+8875 <cjk>
	0xD1: [`\u887D`].string() // U+887D <cjk>
	0xD2: [`\u88B5`].string() // U+88B5 <cjk>
	0xD3: [`\u8872`].string() // U+8872 <cjk>
	0xD4: [`\u8882`].string() // U+8882 <cjk>
	0xD5: [`\u8897`].string() // U+8897 <cjk>
	0xD6: [`\u8892`].string() // U+8892 <cjk>
	0xD7: [`\u88AE`].string() // U+88AE <cjk>
	0xD8: [`\u8899`].string() // U+8899 <cjk>
	0xD9: [`\u88A2`].string() // U+88A2 <cjk>
	0xDA: [`\u888D`].string() // U+888D <cjk>
	0xDB: [`\u88A4`].string() // U+88A4 <cjk>
	0xDC: [`\u88B0`].string() // U+88B0 <cjk>
	0xDD: [`\u88BF`].string() // U+88BF <cjk>
	0xDE: [`\u88B1`].string() // U+88B1 <cjk>
	0xDF: [`\u88C3`].string() // U+88C3 <cjk>
	0xE0: [`\u88C4`].string() // U+88C4 <cjk>
	0xE1: [`\u88D4`].string() // U+88D4 <cjk>
	0xE2: [`\u88D8`].string() // U+88D8 <cjk>
	0xE3: [`\u88D9`].string() // U+88D9 <cjk>
	0xE4: [`\u88DD`].string() // U+88DD <cjk>
	0xE5: [`\u88F9`].string() // U+88F9 <cjk>
	0xE6: [`\u8902`].string() // U+8902 <cjk>
	0xE7: [`\u88FC`].string() // U+88FC <cjk>
	0xE8: [`\u88F4`].string() // U+88F4 <cjk>
	0xE9: [`\u88E8`].string() // U+88E8 <cjk>
	0xEA: [`\u88F2`].string() // U+88F2 <cjk>
	0xEB: [`\u8904`].string() // U+8904 <cjk>
	0xEC: [`\u890C`].string() // U+890C <cjk>
	0xED: [`\u890A`].string() // U+890A <cjk>
	0xEE: [`\u8913`].string() // U+8913 <cjk>
	0xEF: [`\u8943`].string() // U+8943 <cjk>
	0xF0: [`\u891E`].string() // U+891E <cjk>
	0xF1: [`\u8925`].string() // U+8925 <cjk>
	0xF2: [`\u892A`].string() // U+892A <cjk>
	0xF3: [`\u892B`].string() // U+892B <cjk>
	0xF4: [`\u8941`].string() // U+8941 <cjk>
	0xF5: [`\u8944`].string() // U+8944 <cjk>
	0xF6: [`\u893B`].string() // U+893B <cjk>
	0xF7: [`\u8936`].string() // U+8936 <cjk>
	0xF8: [`\u8938`].string() // U+8938 <cjk>
	0xF9: [`\u894C`].string() // U+894C <cjk>
	0xFA: [`\u891D`].string() // U+891D <cjk>
	0xFB: [`\u8960`].string() // U+8960 <cjk>
	0xFC: [`\u895E`].string() // U+895E <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xfc = {
	0x40: [`\u9A31`].string() // U+9A31 <cjk>
	0x41: [`\u9A36`].string() // U+9A36 <cjk>
	0x42: [`\u9A44`].string() // U+9A44 <cjk>
	0x43: [`\u9A4C`].string() // U+9A4C <cjk>
	0x44: [`\u9A58`].string() // U+9A58 <cjk>
	0x45: [`\u4BC2`].string() // U+4BC2 <cjk>
	0x46: [`\u9AAF`].string() // U+9AAF <cjk>
	0x47: [`\u4BCA`].string() // U+4BCA <cjk>
	0x48: [`\u9AB7`].string() // U+9AB7 <cjk>
	0x49: [`\u4BD2`].string() // U+4BD2 <cjk>
	0x4A: [`\u9AB9`].string() // U+9AB9 <cjk>
	0x4B: utf32_to_str(0x29A72) // U+29A72 <cjk>
	0x4C: [`\u9AC6`].string() // U+9AC6 <cjk>
	0x4D: [`\u9AD0`].string() // U+9AD0 <cjk>
	0x4E: [`\u9AD2`].string() // U+9AD2 <cjk>
	0x4F: [`\u9AD5`].string() // U+9AD5 <cjk>
	0x50: [`\u4BE8`].string() // U+4BE8 <cjk>
	0x51: [`\u9ADC`].string() // U+9ADC <cjk>
	0x52: [`\u9AE0`].string() // U+9AE0 <cjk>
	0x53: [`\u9AE5`].string() // U+9AE5 <cjk>
	0x54: [`\u9AE9`].string() // U+9AE9 <cjk>
	0x55: [`\u9B03`].string() // U+9B03 <cjk>
	0x56: [`\u9B0C`].string() // U+9B0C <cjk>
	0x57: [`\u9B10`].string() // U+9B10 <cjk>
	0x58: [`\u9B12`].string() // U+9B12 <cjk>
	0x59: [`\u9B16`].string() // U+9B16 <cjk>
	0x5A: [`\u9B1C`].string() // U+9B1C <cjk>
	0x5B: [`\u9B2B`].string() // U+9B2B <cjk>
	0x5C: [`\u9B33`].string() // U+9B33 <cjk>
	0x5D: [`\u9B3D`].string() // U+9B3D <cjk>
	0x5E: [`\u4C20`].string() // U+4C20 <cjk>
	0x5F: [`\u9B4B`].string() // U+9B4B <cjk>
	0x60: [`\u9B63`].string() // U+9B63 <cjk>
	0x61: [`\u9B65`].string() // U+9B65 <cjk>
	0x62: [`\u9B6B`].string() // U+9B6B <cjk>
	0x63: [`\u9B6C`].string() // U+9B6C <cjk>
	0x64: [`\u9B73`].string() // U+9B73 <cjk>
	0x65: [`\u9B76`].string() // U+9B76 <cjk>
	0x66: [`\u9B77`].string() // U+9B77 <cjk>
	0x67: [`\u9BA6`].string() // U+9BA6 <cjk>
	0x68: [`\u9BAC`].string() // U+9BAC <cjk>
	0x69: [`\u9BB1`].string() // U+9BB1 <cjk>
	0x6A: utf32_to_str(0x29DDB) // U+29DDB <cjk>
	0x6B: utf32_to_str(0x29E3D) // U+29E3D <cjk>
	0x6C: [`\u9BB2`].string() // U+9BB2 <cjk>
	0x6D: [`\u9BB8`].string() // U+9BB8 <cjk>
	0x6E: [`\u9BBE`].string() // U+9BBE <cjk>
	0x6F: [`\u9BC7`].string() // U+9BC7 <cjk>
	0x70: [`\u9BF3`].string() // U+9BF3 <cjk>
	0x71: [`\u9BD8`].string() // U+9BD8 <cjk>
	0x72: [`\u9BDD`].string() // U+9BDD <cjk>
	0x73: [`\u9BE7`].string() // U+9BE7 <cjk>
	0x74: [`\u9BEA`].string() // U+9BEA <cjk>
	0x75: [`\u9BEB`].string() // U+9BEB <cjk>
	0x76: [`\u9BEF`].string() // U+9BEF <cjk>
	0x77: [`\u9BEE`].string() // U+9BEE <cjk>
	0x78: utf32_to_str(0x29E15) // U+29E15 <cjk>
	0x79: [`\u9BFA`].string() // U+9BFA <cjk>
	0x7A: utf32_to_str(0x29E8A) // U+29E8A <cjk>
	0x7B: [`\u9BF7`].string() // U+9BF7 <cjk>
	0x7C: utf32_to_str(0x29E49) // U+29E49 <cjk>
	0x7D: [`\u9C16`].string() // U+9C16 <cjk>
	0x7E: [`\u9C18`].string() // U+9C18 <cjk>
	0x80: [`\u9C19`].string() // U+9C19 <cjk>
	0x81: [`\u9C1A`].string() // U+9C1A <cjk>
	0x82: [`\u9C1D`].string() // U+9C1D <cjk>
	0x83: [`\u9C22`].string() // U+9C22 <cjk>
	0x84: [`\u9C27`].string() // U+9C27 <cjk>
	0x85: [`\u9C29`].string() // U+9C29 <cjk>
	0x86: [`\u9C2A`].string() // U+9C2A <cjk>
	0x87: utf32_to_str(0x29EC4) // U+29EC4 <cjk>
	0x88: [`\u9C31`].string() // U+9C31 <cjk>
	0x89: [`\u9C36`].string() // U+9C36 <cjk>
	0x8A: [`\u9C37`].string() // U+9C37 <cjk>
	0x8B: [`\u9C45`].string() // U+9C45 <cjk>
	0x8C: [`\u9C5C`].string() // U+9C5C <cjk>
	0x8D: utf32_to_str(0x29EE9) // U+29EE9 <cjk>
	0x8E: [`\u9C49`].string() // U+9C49 <cjk>
	0x8F: [`\u9C4A`].string() // U+9C4A <cjk>
	0x90: utf32_to_str(0x29EDB) // U+29EDB <cjk>
	0x91: [`\u9C54`].string() // U+9C54 <cjk>
	0x92: [`\u9C58`].string() // U+9C58 <cjk>
	0x93: [`\u9C5B`].string() // U+9C5B <cjk>
	0x94: [`\u9C5D`].string() // U+9C5D <cjk>
	0x95: [`\u9C5F`].string() // U+9C5F <cjk>
	0x96: [`\u9C69`].string() // U+9C69 <cjk>
	0x97: [`\u9C6A`].string() // U+9C6A <cjk>
	0x98: [`\u9C6B`].string() // U+9C6B <cjk>
	0x99: [`\u9C6D`].string() // U+9C6D <cjk>
	0x9A: [`\u9C6E`].string() // U+9C6E <cjk>
	0x9B: [`\u9C70`].string() // U+9C70 <cjk>
	0x9C: [`\u9C72`].string() // U+9C72 <cjk>
	0x9D: [`\u9C75`].string() // U+9C75 <cjk>
	0x9E: [`\u9C7A`].string() // U+9C7A <cjk>
	0x9F: [`\u9CE6`].string() // U+9CE6 <cjk>
	0xA0: [`\u9CF2`].string() // U+9CF2 <cjk>
	0xA1: [`\u9D0B`].string() // U+9D0B <cjk>
	0xA2: [`\u9D02`].string() // U+9D02 <cjk>
	0xA3: utf32_to_str(0x29FCE) // U+29FCE <cjk>
	0xA4: [`\u9D11`].string() // U+9D11 <cjk>
	0xA5: [`\u9D17`].string() // U+9D17 <cjk>
	0xA6: [`\u9D18`].string() // U+9D18 <cjk>
	0xA7: utf32_to_str(0x2A02F) // U+2A02F <cjk>
	0xA8: [`\u4CC4`].string() // U+4CC4 <cjk>
	0xA9: utf32_to_str(0x2A01A) // U+2A01A <cjk>
	0xAA: [`\u9D32`].string() // U+9D32 <cjk>
	0xAB: [`\u4CD1`].string() // U+4CD1 <cjk>
	0xAC: [`\u9D42`].string() // U+9D42 <cjk>
	0xAD: [`\u9D4A`].string() // U+9D4A <cjk>
	0xAE: [`\u9D5F`].string() // U+9D5F <cjk>
	0xAF: [`\u9D62`].string() // U+9D62 <cjk>
	0xB0: utf32_to_str(0x2A0F9) // U+2A0F9 <cjk>
	0xB1: [`\u9D69`].string() // U+9D69 <cjk>
	0xB2: [`\u9D6B`].string() // U+9D6B <cjk>
	0xB3: utf32_to_str(0x2A082) // U+2A082 <cjk>
	0xB4: [`\u9D73`].string() // U+9D73 <cjk>
	0xB5: [`\u9D76`].string() // U+9D76 <cjk>
	0xB6: [`\u9D77`].string() // U+9D77 <cjk>
	0xB7: [`\u9D7E`].string() // U+9D7E <cjk>
	0xB8: [`\u9D84`].string() // U+9D84 <cjk>
	0xB9: [`\u9D8D`].string() // U+9D8D <cjk>
	0xBA: [`\u9D99`].string() // U+9D99 <cjk>
	0xBB: [`\u9DA1`].string() // U+9DA1 <cjk>
	0xBC: [`\u9DBF`].string() // U+9DBF <cjk>
	0xBD: [`\u9DB5`].string() // U+9DB5 <cjk>
	0xBE: [`\u9DB9`].string() // U+9DB9 <cjk>
	0xBF: [`\u9DBD`].string() // U+9DBD <cjk>
	0xC0: [`\u9DC3`].string() // U+9DC3 <cjk>
	0xC1: [`\u9DC7`].string() // U+9DC7 <cjk>
	0xC2: [`\u9DC9`].string() // U+9DC9 <cjk>
	0xC3: [`\u9DD6`].string() // U+9DD6 <cjk>
	0xC4: [`\u9DDA`].string() // U+9DDA <cjk>
	0xC5: [`\u9DDF`].string() // U+9DDF <cjk>
	0xC6: [`\u9DE0`].string() // U+9DE0 <cjk>
	0xC7: [`\u9DE3`].string() // U+9DE3 <cjk>
	0xC8: [`\u9DF4`].string() // U+9DF4 <cjk>
	0xC9: [`\u4D07`].string() // U+4D07 <cjk>
	0xCA: [`\u9E0A`].string() // U+9E0A <cjk>
	0xCB: [`\u9E02`].string() // U+9E02 <cjk>
	0xCC: [`\u9E0D`].string() // U+9E0D <cjk>
	0xCD: [`\u9E19`].string() // U+9E19 <cjk>
	0xCE: [`\u9E1C`].string() // U+9E1C <cjk>
	0xCF: [`\u9E1D`].string() // U+9E1D <cjk>
	0xD0: [`\u9E7B`].string() // U+9E7B <cjk>
	0xD1: utf32_to_str(0x22218) // U+22218 <cjk>
	0xD2: [`\u9E80`].string() // U+9E80 <cjk>
	0xD3: [`\u9E85`].string() // U+9E85 <cjk>
	0xD4: [`\u9E9B`].string() // U+9E9B <cjk>
	0xD5: [`\u9EA8`].string() // U+9EA8 <cjk>
	0xD6: utf32_to_str(0x2A38C) // U+2A38C <cjk>
	0xD7: [`\u9EBD`].string() // U+9EBD <cjk>
	0xD8: utf32_to_str(0x2A437) // U+2A437 <cjk>
	0xD9: [`\u9EDF`].string() // U+9EDF <cjk>
	0xDA: [`\u9EE7`].string() // U+9EE7 <cjk>
	0xDB: [`\u9EEE`].string() // U+9EEE <cjk>
	0xDC: [`\u9EFF`].string() // U+9EFF <cjk>
	0xDD: [`\u9F02`].string() // U+9F02 <cjk>
	0xDE: [`\u4D77`].string() // U+4D77 <cjk>
	0xDF: [`\u9F03`].string() // U+9F03 <cjk>
	0xE0: [`\u9F17`].string() // U+9F17 <cjk>
	0xE1: [`\u9F19`].string() // U+9F19 <cjk>
	0xE2: [`\u9F2F`].string() // U+9F2F <cjk>
	0xE3: [`\u9F37`].string() // U+9F37 <cjk>
	0xE4: [`\u9F3A`].string() // U+9F3A <cjk>
	0xE5: [`\u9F3D`].string() // U+9F3D <cjk>
	0xE6: [`\u9F41`].string() // U+9F41 <cjk>
	0xE7: [`\u9F45`].string() // U+9F45 <cjk>
	0xE8: [`\u9F46`].string() // U+9F46 <cjk>
	0xE9: [`\u9F53`].string() // U+9F53 <cjk>
	0xEA: [`\u9F55`].string() // U+9F55 <cjk>
	0xEB: [`\u9F58`].string() // U+9F58 <cjk>
	0xEC: utf32_to_str(0x2A5F1) // U+2A5F1 <cjk>
	0xED: [`\u9F5D`].string() // U+9F5D <cjk>
	0xEE: utf32_to_str(0x2A602) // U+2A602 <cjk>
	0xEF: [`\u9F69`].string() // U+9F69 <cjk>
	0xF0: utf32_to_str(0x2A61A) // U+2A61A <cjk>
	0xF1: [`\u9F6D`].string() // U+9F6D <cjk>
	0xF2: [`\u9F70`].string() // U+9F70 <cjk>
	0xF3: [`\u9F75`].string() // U+9F75 <cjk>
	0xF4: utf32_to_str(0x2A6B2) // U+2A6B2 <cjk>
}

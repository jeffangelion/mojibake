module mojibake

const jis_x_0213_doublebyte_0xe1 = {
	0x40: [`\u74E0`].string() // U+74E0 <cjk>
	0x41: [`\u74E3`].string() // U+74E3 <cjk>
	0x42: [`\u74E7`].string() // U+74E7 <cjk>
	0x43: [`\u74E9`].string() // U+74E9 <cjk>
	0x44: [`\u74EE`].string() // U+74EE <cjk>
	0x45: [`\u74F2`].string() // U+74F2 <cjk>
	0x46: [`\u74F0`].string() // U+74F0 <cjk>
	0x47: [`\u74F1`].string() // U+74F1 <cjk>
	0x48: [`\u74F8`].string() // U+74F8 <cjk>
	0x49: [`\u74F7`].string() // U+74F7 <cjk>
	0x4A: [`\u7504`].string() // U+7504 <cjk>
	0x4B: [`\u7503`].string() // U+7503 <cjk>
	0x4C: [`\u7505`].string() // U+7505 <cjk>
	0x4D: [`\u750C`].string() // U+750C <cjk>
	0x4E: [`\u750E`].string() // U+750E <cjk>
	0x4F: [`\u750D`].string() // U+750D <cjk>
	0x50: [`\u7515`].string() // U+7515 <cjk>
	0x51: [`\u7513`].string() // U+7513 <cjk>
	0x52: [`\u751E`].string() // U+751E <cjk>
	0x53: [`\u7526`].string() // U+7526 <cjk>
	0x54: [`\u752C`].string() // U+752C <cjk>
	0x55: [`\u753C`].string() // U+753C <cjk>
	0x56: [`\u7544`].string() // U+7544 <cjk>
	0x57: [`\u754D`].string() // U+754D <cjk>
	0x58: [`\u754A`].string() // U+754A <cjk>
	0x59: [`\u7549`].string() // U+7549 <cjk>
	0x5A: [`\u755B`].string() // U+755B <cjk>
	0x5B: [`\u7546`].string() // U+7546 <cjk>
	0x5C: [`\u755A`].string() // U+755A <cjk>
	0x5D: [`\u7569`].string() // U+7569 <cjk>
	0x5E: [`\u7564`].string() // U+7564 <cjk>
	0x5F: [`\u7567`].string() // U+7567 <cjk>
	0x60: [`\u756B`].string() // U+756B <cjk>
	0x61: [`\u756D`].string() // U+756D <cjk>
	0x62: [`\u7578`].string() // U+7578 <cjk>
	0x63: [`\u7576`].string() // U+7576 <cjk>
	0x64: [`\u7586`].string() // U+7586 <cjk>
	0x65: [`\u7587`].string() // U+7587 <cjk>
	0x66: [`\u7574`].string() // U+7574 <cjk>
	0x67: [`\u758A`].string() // U+758A <cjk>
	0x68: [`\u7589`].string() // U+7589 <cjk>
	0x69: [`\u7582`].string() // U+7582 <cjk>
	0x6A: [`\u7594`].string() // U+7594 <cjk>
	0x6B: [`\u759A`].string() // U+759A <cjk>
	0x6C: [`\u759D`].string() // U+759D <cjk>
	0x6D: [`\u75A5`].string() // U+75A5 <cjk>
	0x6E: [`\u75A3`].string() // U+75A3 <cjk>
	0x6F: [`\u75C2`].string() // U+75C2 <cjk>
	0x70: [`\u75B3`].string() // U+75B3 <cjk>
	0x71: [`\u75C3`].string() // U+75C3 <cjk>
	0x72: [`\u75B5`].string() // U+75B5 <cjk>
	0x73: [`\u75BD`].string() // U+75BD <cjk>
	0x74: [`\u75B8`].string() // U+75B8 <cjk>
	0x75: [`\u75BC`].string() // U+75BC <cjk>
	0x76: [`\u75B1`].string() // U+75B1 <cjk>
	0x77: [`\u75CD`].string() // U+75CD <cjk>
	0x78: [`\u75CA`].string() // U+75CA <cjk>
	0x79: [`\u75D2`].string() // U+75D2 <cjk>
	0x7A: [`\u75D9`].string() // U+75D9 <cjk>
	0x7B: [`\u75E3`].string() // U+75E3 <cjk>
	0x7C: [`\u75DE`].string() // U+75DE <cjk>
	0x7D: [`\u75FE`].string() // U+75FE <cjk>
	0x7E: [`\u75FF`].string() // U+75FF <cjk>
	0x80: [`\u75FC`].string() // U+75FC <cjk>
	0x81: [`\u7601`].string() // U+7601 <cjk>
	0x82: [`\u75F0`].string() // U+75F0 <cjk>
	0x83: [`\u75FA`].string() // U+75FA <cjk>
	0x84: [`\u75F2`].string() // U+75F2 <cjk>
	0x85: [`\u75F3`].string() // U+75F3 <cjk>
	0x86: [`\u760B`].string() // U+760B <cjk>
	0x87: [`\u760D`].string() // U+760D <cjk>
	0x88: [`\u7609`].string() // U+7609 <cjk>
	0x89: [`\u761F`].string() // U+761F <cjk>
	0x8A: [`\u7627`].string() // U+7627 <cjk>
	0x8B: [`\u7620`].string() // U+7620 <cjk>
	0x8C: [`\u7621`].string() // U+7621 <cjk>
	0x8D: [`\u7622`].string() // U+7622 <cjk>
	0x8E: [`\u7624`].string() // U+7624 <cjk>
	0x8F: [`\u7634`].string() // U+7634 <cjk>
	0x90: [`\u7630`].string() // U+7630 <cjk>
	0x91: [`\u763B`].string() // U+763B <cjk>
	0x92: [`\u7647`].string() // U+7647 <cjk>
	0x93: [`\u7648`].string() // U+7648 <cjk>
	0x94: [`\u7646`].string() // U+7646 <cjk>
	0x95: [`\u765C`].string() // U+765C <cjk>
	0x96: [`\u7658`].string() // U+7658 <cjk>
	0x97: [`\u7661`].string() // U+7661 <cjk>
	0x98: [`\u7662`].string() // U+7662 <cjk>
	0x99: [`\u7668`].string() // U+7668 <cjk>
	0x9A: [`\u7669`].string() // U+7669 <cjk>
	0x9B: [`\u766A`].string() // U+766A <cjk>
	0x9C: [`\u7667`].string() // U+7667 <cjk>
	0x9D: [`\u766C`].string() // U+766C <cjk>
	0x9E: [`\u7670`].string() // U+7670 <cjk>
	0x9F: [`\u7672`].string() // U+7672 <cjk>
	0xA0: [`\u7676`].string() // U+7676 <cjk>
	0xA1: [`\u7678`].string() // U+7678 <cjk>
	0xA2: [`\u767C`].string() // U+767C <cjk>
	0xA3: [`\u7680`].string() // U+7680 <cjk>
	0xA4: [`\u7683`].string() // U+7683 <cjk>
	0xA5: [`\u7688`].string() // U+7688 <cjk>
	0xA6: [`\u768B`].string() // U+768B <cjk>
	0xA7: [`\u768E`].string() // U+768E <cjk>
	0xA8: [`\u7696`].string() // U+7696 <cjk>
	0xA9: [`\u7693`].string() // U+7693 <cjk>
	0xAA: [`\u7699`].string() // U+7699 <cjk>
	0xAB: [`\u769A`].string() // U+769A <cjk>
	0xAC: [`\u76B0`].string() // U+76B0 <cjk>
	0xAD: [`\u76B4`].string() // U+76B4 <cjk>
	0xAE: [`\u76B8`].string() // U+76B8 <cjk>
	0xAF: [`\u76B9`].string() // U+76B9 <cjk>
	0xB0: [`\u76BA`].string() // U+76BA <cjk>
	0xB1: [`\u76C2`].string() // U+76C2 <cjk>
	0xB2: [`\u76CD`].string() // U+76CD <cjk>
	0xB3: [`\u76D6`].string() // U+76D6 <cjk>
	0xB4: [`\u76D2`].string() // U+76D2 <cjk>
	0xB5: [`\u76DE`].string() // U+76DE <cjk>
	0xB6: [`\u76E1`].string() // U+76E1 <cjk>
	0xB7: [`\u76E5`].string() // U+76E5 <cjk>
	0xB8: [`\u76E7`].string() // U+76E7 <cjk>
	0xB9: [`\u76EA`].string() // U+76EA <cjk>
	0xBA: [`\u862F`].string() // U+862F <cjk>
	0xBB: [`\u76FB`].string() // U+76FB <cjk>
	0xBC: [`\u7708`].string() // U+7708 <cjk>
	0xBD: [`\u7707`].string() // U+7707 <cjk>
	0xBE: [`\u7704`].string() // U+7704 <cjk>
	0xBF: [`\u7729`].string() // U+7729 <cjk>
	0xC0: [`\u7724`].string() // U+7724 <cjk>
	0xC1: [`\u771E`].string() // U+771E <cjk>
	0xC2: [`\u7725`].string() // U+7725 <cjk>
	0xC3: [`\u7726`].string() // U+7726 <cjk>
	0xC4: [`\u771B`].string() // U+771B <cjk>
	0xC5: [`\u7737`].string() // U+7737 <cjk>
	0xC6: [`\u7738`].string() // U+7738 <cjk>
	0xC7: [`\u7747`].string() // U+7747 <cjk>
	0xC8: [`\u775A`].string() // U+775A <cjk>
	0xC9: [`\u7768`].string() // U+7768 <cjk>
	0xCA: [`\u776B`].string() // U+776B <cjk>
	0xCB: [`\u775B`].string() // U+775B <cjk>
	0xCC: [`\u7765`].string() // U+7765 <cjk>
	0xCD: [`\u777F`].string() // U+777F <cjk>
	0xCE: [`\u777E`].string() // U+777E <cjk>
	0xCF: [`\u7779`].string() // U+7779 <cjk>
	0xD0: [`\u778E`].string() // U+778E <cjk>
	0xD1: [`\u778B`].string() // U+778B <cjk>
	0xD2: [`\u7791`].string() // U+7791 <cjk>
	0xD3: [`\u77A0`].string() // U+77A0 <cjk>
	0xD4: [`\u779E`].string() // U+779E <cjk>
	0xD5: [`\u77B0`].string() // U+77B0 <cjk>
	0xD6: [`\u77B6`].string() // U+77B6 <cjk>
	0xD7: [`\u77B9`].string() // U+77B9 <cjk>
	0xD8: [`\u77BF`].string() // U+77BF <cjk>
	0xD9: [`\u77BC`].string() // U+77BC <cjk>
	0xDA: [`\u77BD`].string() // U+77BD <cjk>
	0xDB: [`\u77BB`].string() // U+77BB <cjk>
	0xDC: [`\u77C7`].string() // U+77C7 <cjk>
	0xDD: [`\u77CD`].string() // U+77CD <cjk>
	0xDE: [`\u77D7`].string() // U+77D7 <cjk>
	0xDF: [`\u77DA`].string() // U+77DA <cjk>
	0xE0: [`\u77DC`].string() // U+77DC <cjk>
	0xE1: [`\u77E3`].string() // U+77E3 <cjk>
	0xE2: [`\u77EE`].string() // U+77EE <cjk>
	0xE3: [`\u77FC`].string() // U+77FC <cjk>
	0xE4: [`\u780C`].string() // U+780C <cjk>
	0xE5: [`\u7812`].string() // U+7812 <cjk>
	0xE6: [`\u7926`].string() // U+7926 <cjk>
	0xE7: [`\u7820`].string() // U+7820 <cjk>
	0xE8: [`\u792A`].string() // U+792A <cjk>
	0xE9: [`\u7845`].string() // U+7845 <cjk>
	0xEA: [`\u788E`].string() // U+788E <cjk>
	0xEB: [`\u7874`].string() // U+7874 <cjk>
	0xEC: [`\u7886`].string() // U+7886 <cjk>
	0xED: [`\u787C`].string() // U+787C <cjk>
	0xEE: [`\u789A`].string() // U+789A <cjk>
	0xEF: [`\u788C`].string() // U+788C <cjk>
	0xF0: [`\u78A3`].string() // U+78A3 <cjk>
	0xF1: [`\u78B5`].string() // U+78B5 <cjk>
	0xF2: [`\u78AA`].string() // U+78AA <cjk>
	0xF3: [`\u78AF`].string() // U+78AF <cjk>
	0xF4: [`\u78D1`].string() // U+78D1 <cjk>
	0xF5: [`\u78C6`].string() // U+78C6 <cjk>
	0xF6: [`\u78CB`].string() // U+78CB <cjk>
	0xF7: [`\u78D4`].string() // U+78D4 <cjk>
	0xF8: [`\u78BE`].string() // U+78BE <cjk>
	0xF9: [`\u78BC`].string() // U+78BC <cjk>
	0xFA: [`\u78C5`].string() // U+78C5 <cjk>
	0xFB: [`\u78CA`].string() // U+78CA <cjk>
	0xFC: [`\u78EC`].string() // U+78EC <cjk>
}

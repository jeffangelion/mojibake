module mojibake

const jis_x_0213_doublebyte_0x95 = {
	0x40: [`\u9F3B`].string() // U+9F3B <cjk>
	0x41: [`\u67CA`].string() // U+67CA <cjk>
	0x42: [`\u7A17`].string() // U+7A17 <cjk>
	0x43: [`\u5339`].string() // U+5339 <cjk>
	0x44: [`\u758B`].string() // U+758B <cjk>
	0x45: [`\u9AED`].string() // U+9AED <cjk>
	0x46: [`\u5F66`].string() // U+5F66 <cjk>
	0x47: [`\u819D`].string() // U+819D <cjk>
	0x48: [`\u83F1`].string() // U+83F1 <cjk>
	0x49: [`\u8098`].string() // U+8098 <cjk>
	0x4A: [`\u5F3C`].string() // U+5F3C <cjk>
	0x4B: [`\u5FC5`].string() // U+5FC5 <cjk>
	0x4C: [`\u7562`].string() // U+7562 <cjk>
	0x4D: [`\u7B46`].string() // U+7B46 <cjk>
	0x4E: [`\u903C`].string() // U+903C <cjk>
	0x4F: [`\u6867`].string() // U+6867 <cjk>
	0x50: [`\u59EB`].string() // U+59EB <cjk>
	0x51: [`\u5A9B`].string() // U+5A9B <cjk>
	0x52: [`\u7D10`].string() // U+7D10 <cjk>
	0x53: [`\u767E`].string() // U+767E <cjk>
	0x54: [`\u8B2C`].string() // U+8B2C <cjk>
	0x55: [`\u4FF5`].string() // U+4FF5 <cjk>
	0x56: [`\u5F6A`].string() // U+5F6A <cjk>
	0x57: [`\u6A19`].string() // U+6A19 <cjk>
	0x58: [`\u6C37`].string() // U+6C37 <cjk>
	0x59: [`\u6F02`].string() // U+6F02 <cjk>
	0x5A: [`\u74E2`].string() // U+74E2 <cjk>
	0x5B: [`\u7968`].string() // U+7968 <cjk>
	0x5C: [`\u8868`].string() // U+8868 <cjk>
	0x5D: [`\u8A55`].string() // U+8A55 <cjk>
	0x5E: [`\u8C79`].string() // U+8C79 <cjk>
	0x5F: [`\u5EDF`].string() // U+5EDF <cjk>
	0x60: [`\u63CF`].string() // U+63CF <cjk>
	0x61: [`\u75C5`].string() // U+75C5 <cjk>
	0x62: [`\u79D2`].string() // U+79D2 <cjk>
	0x63: [`\u82D7`].string() // U+82D7 <cjk>
	0x64: [`\u9328`].string() // U+9328 <cjk>
	0x65: [`\u92F2`].string() // U+92F2 <cjk>
	0x66: [`\u849C`].string() // U+849C <cjk>
	0x67: [`\u86ED`].string() // U+86ED <cjk>
	0x68: [`\u9C2D`].string() // U+9C2D <cjk>
	0x69: [`\u54C1`].string() // U+54C1 <cjk>
	0x6A: [`\u5F6C`].string() // U+5F6C <cjk>
	0x6B: [`\u658C`].string() // U+658C <cjk>
	0x6C: [`\u6D5C`].string() // U+6D5C <cjk>
	0x6D: [`\u7015`].string() // U+7015 <cjk>
	0x6E: [`\u8CA7`].string() // U+8CA7 <cjk>
	0x6F: [`\u8CD3`].string() // U+8CD3 <cjk>
	0x70: [`\u983B`].string() // U+983B <cjk>
	0x71: [`\u654F`].string() // U+654F <cjk>
	0x72: [`\u74F6`].string() // U+74F6 <cjk>
	0x73: [`\u4E0D`].string() // U+4E0D <cjk>
	0x74: [`\u4ED8`].string() // U+4ED8 <cjk>
	0x75: [`\u57E0`].string() // U+57E0 <cjk>
	0x76: [`\u592B`].string() // U+592B <cjk>
	0x77: [`\u5A66`].string() // U+5A66 <cjk>
	0x78: [`\u5BCC`].string() // U+5BCC <cjk>
	0x79: [`\u51A8`].string() // U+51A8 <cjk>
	0x7A: [`\u5E03`].string() // U+5E03 <cjk>
	0x7B: [`\u5E9C`].string() // U+5E9C <cjk>
	0x7C: [`\u6016`].string() // U+6016 <cjk>
	0x7D: [`\u6276`].string() // U+6276 <cjk>
	0x7E: [`\u6577`].string() // U+6577 <cjk>
	0x80: [`\u65A7`].string() // U+65A7 <cjk>
	0x81: [`\u666E`].string() // U+666E <cjk>
	0x82: [`\u6D6E`].string() // U+6D6E <cjk>
	0x83: [`\u7236`].string() // U+7236 <cjk>
	0x84: [`\u7B26`].string() // U+7B26 <cjk>
	0x85: [`\u8150`].string() // U+8150 <cjk>
	0x86: [`\u819A`].string() // U+819A <cjk>
	0x87: [`\u8299`].string() // U+8299 <cjk>
	0x88: [`\u8B5C`].string() // U+8B5C <cjk>
	0x89: [`\u8CA0`].string() // U+8CA0 <cjk>
	0x8A: [`\u8CE6`].string() // U+8CE6 <cjk>
	0x8B: [`\u8D74`].string() // U+8D74 <cjk>
	0x8C: [`\u961C`].string() // U+961C <cjk>
	0x8D: [`\u9644`].string() // U+9644 <cjk>
	0x8E: [`\u4FAE`].string() // U+4FAE <cjk>
	0x8F: [`\u64AB`].string() // U+64AB <cjk>
	0x90: [`\u6B66`].string() // U+6B66 <cjk>
	0x91: [`\u821E`].string() // U+821E <cjk>
	0x92: [`\u8461`].string() // U+8461 <cjk>
	0x93: [`\u856A`].string() // U+856A <cjk>
	0x94: [`\u90E8`].string() // U+90E8 <cjk>
	0x95: [`\u5C01`].string() // U+5C01 <cjk>
	0x96: [`\u6953`].string() // U+6953 <cjk>
	0x97: [`\u98A8`].string() // U+98A8 <cjk>
	0x98: [`\u847A`].string() // U+847A <cjk>
	0x99: [`\u8557`].string() // U+8557 <cjk>
	0x9A: [`\u4F0F`].string() // U+4F0F <cjk>
	0x9B: [`\u526F`].string() // U+526F <cjk>
	0x9C: [`\u5FA9`].string() // U+5FA9 <cjk>
	0x9D: [`\u5E45`].string() // U+5E45 <cjk>
	0x9E: [`\u670D`].string() // U+670D <cjk>
	0x9F: [`\u798F`].string() // U+798F <cjk>
	0xA0: [`\u8179`].string() // U+8179 <cjk>
	0xA1: [`\u8907`].string() // U+8907 <cjk>
	0xA2: [`\u8986`].string() // U+8986 <cjk>
	0xA3: [`\u6DF5`].string() // U+6DF5 <cjk>
	0xA4: [`\u5F17`].string() // U+5F17 <cjk>
	0xA5: [`\u6255`].string() // U+6255 <cjk>
	0xA6: [`\u6CB8`].string() // U+6CB8 <cjk>
	0xA7: [`\u4ECF`].string() // U+4ECF <cjk>
	0xA8: [`\u7269`].string() // U+7269 <cjk>
	0xA9: [`\u9B92`].string() // U+9B92 <cjk>
	0xAA: [`\u5206`].string() // U+5206 <cjk>
	0xAB: [`\u543B`].string() // U+543B <cjk>
	0xAC: [`\u5674`].string() // U+5674 <cjk>
	0xAD: [`\u58B3`].string() // U+58B3 <cjk>
	0xAE: [`\u61A4`].string() // U+61A4 <cjk>
	0xAF: [`\u626E`].string() // U+626E <cjk>
	0xB0: [`\u711A`].string() // U+711A <cjk>
	0xB1: [`\u596E`].string() // U+596E <cjk>
	0xB2: [`\u7C89`].string() // U+7C89 <cjk>
	0xB3: [`\u7CDE`].string() // U+7CDE <cjk>
	0xB4: [`\u7D1B`].string() // U+7D1B <cjk>
	0xB5: [`\u96F0`].string() // U+96F0 <cjk>
	0xB6: [`\u6587`].string() // U+6587 <cjk>
	0xB7: [`\u805E`].string() // U+805E <cjk>
	0xB8: [`\u4E19`].string() // U+4E19 <cjk>
	0xB9: [`\u4F75`].string() // U+4F75 <cjk>
	0xBA: [`\u5175`].string() // U+5175 <cjk>
	0xBB: [`\u5840`].string() // U+5840 <cjk>
	0xBC: [`\u5E63`].string() // U+5E63 <cjk>
	0xBD: [`\u5E73`].string() // U+5E73 <cjk>
	0xBE: [`\u5F0A`].string() // U+5F0A <cjk>
	0xBF: [`\u67C4`].string() // U+67C4 <cjk>
	0xC0: [`\u4E26`].string() // U+4E26 <cjk>
	0xC1: [`\u853D`].string() // U+853D <cjk>
	0xC2: [`\u9589`].string() // U+9589 <cjk>
	0xC3: [`\u965B`].string() // U+965B <cjk>
	0xC4: [`\u7C73`].string() // U+7C73 <cjk>
	0xC5: [`\u9801`].string() // U+9801 <cjk>
	0xC6: [`\u50FB`].string() // U+50FB <cjk>
	0xC7: [`\u58C1`].string() // U+58C1 <cjk>
	0xC8: [`\u7656`].string() // U+7656 <cjk>
	0xC9: [`\u78A7`].string() // U+78A7 <cjk>
	0xCA: [`\u5225`].string() // U+5225 <cjk>
	0xCB: [`\u77A5`].string() // U+77A5 <cjk>
	0xCC: [`\u8511`].string() // U+8511 <cjk>
	0xCD: [`\u7B86`].string() // U+7B86 <cjk>
	0xCE: [`\u504F`].string() // U+504F <cjk>
	0xCF: [`\u5909`].string() // U+5909 <cjk>
	0xD0: [`\u7247`].string() // U+7247 <cjk>
	0xD1: [`\u7BC7`].string() // U+7BC7 <cjk>
	0xD2: [`\u7DE8`].string() // U+7DE8 <cjk>
	0xD3: [`\u8FBA`].string() // U+8FBA <cjk>
	0xD4: [`\u8FD4`].string() // U+8FD4 <cjk>
	0xD5: [`\u904D`].string() // U+904D <cjk>
	0xD6: [`\u4FBF`].string() // U+4FBF <cjk>
	0xD7: [`\u52C9`].string() // U+52C9 <cjk>
	0xD8: [`\u5A29`].string() // U+5A29 <cjk>
	0xD9: [`\u5F01`].string() // U+5F01 <cjk>
	0xDA: [`\u97AD`].string() // U+97AD <cjk>
	0xDB: [`\u4FDD`].string() // U+4FDD <cjk>
	0xDC: [`\u8217`].string() // U+8217 <cjk>
	0xDD: [`\u92EA`].string() // U+92EA <cjk>
	0xDE: [`\u5703`].string() // U+5703 <cjk>
	0xDF: [`\u6355`].string() // U+6355 <cjk>
	0xE0: [`\u6B69`].string() // U+6B69 <cjk>
	0xE1: [`\u752B`].string() // U+752B <cjk>
	0xE2: [`\u88DC`].string() // U+88DC <cjk>
	0xE3: [`\u8F14`].string() // U+8F14 <cjk>
	0xE4: [`\u7A42`].string() // U+7A42 <cjk>
	0xE5: [`\u52DF`].string() // U+52DF <cjk>
	0xE6: [`\u5893`].string() // U+5893 <cjk>
	0xE7: [`\u6155`].string() // U+6155 <cjk>
	0xE8: [`\u620A`].string() // U+620A <cjk>
	0xE9: [`\u66AE`].string() // U+66AE <cjk>
	0xEA: [`\u6BCD`].string() // U+6BCD <cjk>
	0xEB: [`\u7C3F`].string() // U+7C3F <cjk>
	0xEC: [`\u83E9`].string() // U+83E9 <cjk>
	0xED: [`\u5023`].string() // U+5023 <cjk>
	0xEE: [`\u4FF8`].string() // U+4FF8 <cjk>
	0xEF: [`\u5305`].string() // U+5305 <cjk>
	0xF0: [`\u5446`].string() // U+5446 <cjk>
	0xF1: [`\u5831`].string() // U+5831 <cjk>
	0xF2: [`\u5949`].string() // U+5949 <cjk>
	0xF3: [`\u5B9D`].string() // U+5B9D <cjk>
	0xF4: [`\u5CF0`].string() // U+5CF0 <cjk>
	0xF5: [`\u5CEF`].string() // U+5CEF <cjk>
	0xF6: [`\u5D29`].string() // U+5D29 <cjk>
	0xF7: [`\u5E96`].string() // U+5E96 <cjk>
	0xF8: [`\u62B1`].string() // U+62B1 <cjk>
	0xF9: [`\u6367`].string() // U+6367 <cjk>
	0xFA: [`\u653E`].string() // U+653E <cjk>
	0xFB: [`\u65B9`].string() // U+65B9 <cjk>
	0xFC: [`\u670B`].string() // U+670B <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xf7 = {
	0x40: [`\u7A38`].string() // U+7A38 <cjk>
	0x41: [`\u7A47`].string() // U+7A47 <cjk>
	0x42: [`\u7A4C`].string() // U+7A4C <cjk>
	0x43: [`\u7A56`].string() // U+7A56 <cjk>
	0x44: [`\u7A59`].string() // U+7A59 <cjk>
	0x45: [`\u7A5C`].string() // U+7A5C <cjk>
	0x46: [`\u7A5F`].string() // U+7A5F <cjk>
	0x47: [`\u7A60`].string() // U+7A60 <cjk>
	0x48: [`\u7A67`].string() // U+7A67 <cjk>
	0x49: [`\u7A6A`].string() // U+7A6A <cjk>
	0x4A: [`\u7A75`].string() // U+7A75 <cjk>
	0x4B: [`\u7A78`].string() // U+7A78 <cjk>
	0x4C: [`\u7A82`].string() // U+7A82 <cjk>
	0x4D: [`\u7A8A`].string() // U+7A8A <cjk>
	0x4E: [`\u7A90`].string() // U+7A90 <cjk>
	0x4F: [`\u7AA3`].string() // U+7AA3 <cjk>
	0x50: [`\u7AAC`].string() // U+7AAC <cjk>
	0x51: utf32_to_str(0x259D4) // U+259D4 <cjk>
	0x52: [`\u41B4`].string() // U+41B4 <cjk>
	0x53: [`\u7AB9`].string() // U+7AB9 <cjk>
	0x54: [`\u7ABC`].string() // U+7ABC <cjk>
	0x55: [`\u7ABE`].string() // U+7ABE <cjk>
	0x56: [`\u41BF`].string() // U+41BF <cjk>
	0x57: [`\u7ACC`].string() // U+7ACC <cjk>
	0x58: [`\u7AD1`].string() // U+7AD1 <cjk>
	0x59: [`\u7AE7`].string() // U+7AE7 <cjk>
	0x5A: [`\u7AE8`].string() // U+7AE8 <cjk>
	0x5B: [`\u7AF4`].string() // U+7AF4 <cjk>
	0x5C: utf32_to_str(0x25AE4) // U+25AE4 <cjk>
	0x5D: utf32_to_str(0x25AE3) // U+25AE3 <cjk>
	0x5E: [`\u7B07`].string() // U+7B07 <cjk>
	0x5F: utf32_to_str(0x25AF1) // U+25AF1 <cjk>
	0x60: [`\u7B3D`].string() // U+7B3D <cjk>
	0x61: [`\u7B27`].string() // U+7B27 <cjk>
	0x62: [`\u7B2A`].string() // U+7B2A <cjk>
	0x63: [`\u7B2E`].string() // U+7B2E <cjk>
	0x64: [`\u7B2F`].string() // U+7B2F <cjk>
	0x65: [`\u7B31`].string() // U+7B31 <cjk>
	0x66: [`\u41E6`].string() // U+41E6 <cjk>
	0x67: [`\u41F3`].string() // U+41F3 <cjk>
	0x68: [`\u7B7F`].string() // U+7B7F <cjk>
	0x69: [`\u7B41`].string() // U+7B41 <cjk>
	0x6A: [`\u41EE`].string() // U+41EE <cjk>
	0x6B: [`\u7B55`].string() // U+7B55 <cjk>
	0x6C: [`\u7B79`].string() // U+7B79 <cjk>
	0x6D: [`\u7B64`].string() // U+7B64 <cjk>
	0x6E: [`\u7B66`].string() // U+7B66 <cjk>
	0x6F: [`\u7B69`].string() // U+7B69 <cjk>
	0x70: [`\u7B73`].string() // U+7B73 <cjk>
	0x71: utf32_to_str(0x25BB2) // U+25BB2 <cjk>
	0x72: [`\u4207`].string() // U+4207 <cjk>
	0x73: [`\u7B90`].string() // U+7B90 <cjk>
	0x74: [`\u7B91`].string() // U+7B91 <cjk>
	0x75: [`\u7B9B`].string() // U+7B9B <cjk>
	0x76: [`\u420E`].string() // U+420E <cjk>
	0x77: [`\u7BAF`].string() // U+7BAF <cjk>
	0x78: [`\u7BB5`].string() // U+7BB5 <cjk>
	0x79: [`\u7BBC`].string() // U+7BBC <cjk>
	0x7A: [`\u7BC5`].string() // U+7BC5 <cjk>
	0x7B: [`\u7BCA`].string() // U+7BCA <cjk>
	0x7C: utf32_to_str(0x25C4B) // U+25C4B <cjk>
	0x7D: utf32_to_str(0x25C64) // U+25C64 <cjk>
	0x7E: [`\u7BD4`].string() // U+7BD4 <cjk>
	0x80: [`\u7BD6`].string() // U+7BD6 <cjk>
	0x81: [`\u7BDA`].string() // U+7BDA <cjk>
	0x82: [`\u7BEA`].string() // U+7BEA <cjk>
	0x83: [`\u7BF0`].string() // U+7BF0 <cjk>
	0x84: [`\u7C03`].string() // U+7C03 <cjk>
	0x85: [`\u7C0B`].string() // U+7C0B <cjk>
	0x86: [`\u7C0E`].string() // U+7C0E <cjk>
	0x87: [`\u7C0F`].string() // U+7C0F <cjk>
	0x88: [`\u7C26`].string() // U+7C26 <cjk>
	0x89: [`\u7C45`].string() // U+7C45 <cjk>
	0x8A: [`\u7C4A`].string() // U+7C4A <cjk>
	0x8B: [`\u7C51`].string() // U+7C51 <cjk>
	0x8C: [`\u7C57`].string() // U+7C57 <cjk>
	0x8D: [`\u7C5E`].string() // U+7C5E <cjk>
	0x8E: [`\u7C61`].string() // U+7C61 <cjk>
	0x8F: [`\u7C69`].string() // U+7C69 <cjk>
	0x90: [`\u7C6E`].string() // U+7C6E <cjk>
	0x91: [`\u7C6F`].string() // U+7C6F <cjk>
	0x92: [`\u7C70`].string() // U+7C70 <cjk>
	0x93: utf32_to_str(0x25E2E) // U+25E2E <cjk>
	0x94: utf32_to_str(0x25E56) // U+25E56 <cjk>
	0x95: utf32_to_str(0x25E65) // U+25E65 <cjk>
	0x96: [`\u7CA6`].string() // U+7CA6 <cjk>
	0x97: utf32_to_str(0x25E62) // U+25E62 <cjk>
	0x98: [`\u7CB6`].string() // U+7CB6 <cjk>
	0x99: [`\u7CB7`].string() // U+7CB7 <cjk>
	0x9A: [`\u7CBF`].string() // U+7CBF <cjk>
	0x9B: utf32_to_str(0x25ED8) // U+25ED8 <cjk>
	0x9C: [`\u7CC4`].string() // U+7CC4 <cjk>
	0x9D: utf32_to_str(0x25EC2) // U+25EC2 <cjk>
	0x9E: [`\u7CC8`].string() // U+7CC8 <cjk>
	0x9F: [`\u7CCD`].string() // U+7CCD <cjk>
	0xA0: utf32_to_str(0x25EE8) // U+25EE8 <cjk>
	0xA1: [`\u7CD7`].string() // U+7CD7 <cjk>
	0xA2: utf32_to_str(0x25F23) // U+25F23 <cjk>
	0xA3: [`\u7CE6`].string() // U+7CE6 <cjk>
	0xA4: [`\u7CEB`].string() // U+7CEB <cjk>
	0xA5: utf32_to_str(0x25F5C) // U+25F5C <cjk>
	0xA6: [`\u7CF5`].string() // U+7CF5 <cjk>
	0xA7: [`\u7D03`].string() // U+7D03 <cjk>
	0xA8: [`\u7D09`].string() // U+7D09 <cjk>
	0xA9: [`\u42C6`].string() // U+42C6 <cjk>
	0xAA: [`\u7D12`].string() // U+7D12 <cjk>
	0xAB: [`\u7D1E`].string() // U+7D1E <cjk>
	0xAC: utf32_to_str(0x25FE0) // U+25FE0 <cjk>
	0xAD: utf32_to_str(0x25FD4) // U+25FD4 <cjk>
	0xAE: [`\u7D3D`].string() // U+7D3D <cjk>
	0xAF: [`\u7D3E`].string() // U+7D3E <cjk>
	0xB0: [`\u7D40`].string() // U+7D40 <cjk>
	0xB1: [`\u7D47`].string() // U+7D47 <cjk>
	0xB2: utf32_to_str(0x2600C) // U+2600C <cjk>
	0xB3: utf32_to_str(0x25FFB) // U+25FFB <cjk>
	0xB4: [`\u42D6`].string() // U+42D6 <cjk>
	0xB5: [`\u7D59`].string() // U+7D59 <cjk>
	0xB6: [`\u7D5A`].string() // U+7D5A <cjk>
	0xB7: [`\u7D6A`].string() // U+7D6A <cjk>
	0xB8: [`\u7D70`].string() // U+7D70 <cjk>
	0xB9: [`\u42DD`].string() // U+42DD <cjk>
	0xBA: [`\u7D7F`].string() // U+7D7F <cjk>
	0xBB: utf32_to_str(0x26017) // U+26017 <cjk>
	0xBC: [`\u7D86`].string() // U+7D86 <cjk>
	0xBD: [`\u7D88`].string() // U+7D88 <cjk>
	0xBE: [`\u7D8C`].string() // U+7D8C <cjk>
	0xBF: [`\u7D97`].string() // U+7D97 <cjk>
	0xC0: utf32_to_str(0x26060) // U+26060 <cjk>
	0xC1: [`\u7D9D`].string() // U+7D9D <cjk>
	0xC2: [`\u7DA7`].string() // U+7DA7 <cjk>
	0xC3: [`\u7DAA`].string() // U+7DAA <cjk>
	0xC4: [`\u7DB6`].string() // U+7DB6 <cjk>
	0xC5: [`\u7DB7`].string() // U+7DB7 <cjk>
	0xC6: [`\u7DC0`].string() // U+7DC0 <cjk>
	0xC7: [`\u7DD7`].string() // U+7DD7 <cjk>
	0xC8: [`\u7DD9`].string() // U+7DD9 <cjk>
	0xC9: [`\u7DE6`].string() // U+7DE6 <cjk>
	0xCA: [`\u7DF1`].string() // U+7DF1 <cjk>
	0xCB: [`\u7DF9`].string() // U+7DF9 <cjk>
	0xCC: [`\u4302`].string() // U+4302 <cjk>
	0xCD: utf32_to_str(0x260ED) // U+260ED <cjk>
	0xCE: [`\uFA58`].string() // U+FA58 CJK COMPATIBILITY IDEOGRAPH-FA58
	0xCF: [`\u7E10`].string() // U+7E10 <cjk>
	0xD0: [`\u7E17`].string() // U+7E17 <cjk>
	0xD1: [`\u7E1D`].string() // U+7E1D <cjk>
	0xD2: [`\u7E20`].string() // U+7E20 <cjk>
	0xD3: [`\u7E27`].string() // U+7E27 <cjk>
	0xD4: [`\u7E2C`].string() // U+7E2C <cjk>
	0xD5: [`\u7E45`].string() // U+7E45 <cjk>
	0xD6: [`\u7E73`].string() // U+7E73 <cjk>
	0xD7: [`\u7E75`].string() // U+7E75 <cjk>
	0xD8: [`\u7E7E`].string() // U+7E7E <cjk>
	0xD9: [`\u7E86`].string() // U+7E86 <cjk>
	0xDA: [`\u7E87`].string() // U+7E87 <cjk>
	0xDB: [`\u432B`].string() // U+432B <cjk>
	0xDC: [`\u7E91`].string() // U+7E91 <cjk>
	0xDD: [`\u7E98`].string() // U+7E98 <cjk>
	0xDE: [`\u7E9A`].string() // U+7E9A <cjk>
	0xDF: [`\u4343`].string() // U+4343 <cjk>
	0xE0: [`\u7F3C`].string() // U+7F3C <cjk>
	0xE1: [`\u7F3B`].string() // U+7F3B <cjk>
	0xE2: [`\u7F3E`].string() // U+7F3E <cjk>
	0xE3: [`\u7F43`].string() // U+7F43 <cjk>
	0xE4: [`\u7F44`].string() // U+7F44 <cjk>
	0xE5: [`\u7F4F`].string() // U+7F4F <cjk>
	0xE6: [`\u34C1`].string() // U+34C1 <cjk>
	0xE7: utf32_to_str(0x26270) // U+26270 <cjk>
	0xE8: [`\u7F52`].string() // U+7F52 <cjk>
	0xE9: utf32_to_str(0x26286) // U+26286 <cjk>
	0xEA: [`\u7F61`].string() // U+7F61 <cjk>
	0xEB: [`\u7F63`].string() // U+7F63 <cjk>
	0xEC: [`\u7F64`].string() // U+7F64 <cjk>
	0xED: [`\u7F6D`].string() // U+7F6D <cjk>
	0xEE: [`\u7F7D`].string() // U+7F7D <cjk>
	0xEF: [`\u7F7E`].string() // U+7F7E <cjk>
	0xF0: utf32_to_str(0x2634C) // U+2634C <cjk>
	0xF1: [`\u7F90`].string() // U+7F90 <cjk>
	0xF2: [`\u517B`].string() // U+517B <cjk>
	0xF3: utf32_to_str(0x23D0E) // U+23D0E <cjk>
	0xF4: [`\u7F96`].string() // U+7F96 <cjk>
	0xF5: [`\u7F9C`].string() // U+7F9C <cjk>
	0xF6: [`\u7FAD`].string() // U+7FAD <cjk>
	0xF7: utf32_to_str(0x26402) // U+26402 <cjk>
	0xF8: [`\u7FC3`].string() // U+7FC3 <cjk>
	0xF9: [`\u7FCF`].string() // U+7FCF <cjk>
	0xFA: [`\u7FE3`].string() // U+7FE3 <cjk>
	0xFB: [`\u7FE5`].string() // U+7FE5 <cjk>
	0xFC: [`\u7FEF`].string() // U+7FEF <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x98 = {
	0x40: [`\u84EE`].string() // U+84EE <cjk>
	0x41: [`\u9023`].string() // U+9023 <cjk>
	0x42: [`\u932C`].string() // U+932C <cjk>
	0x43: [`\u5442`].string() // U+5442 <cjk>
	0x44: [`\u9B6F`].string() // U+9B6F <cjk>
	0x45: [`\u6AD3`].string() // U+6AD3 <cjk>
	0x46: [`\u7089`].string() // U+7089 <cjk>
	0x47: [`\u8CC2`].string() // U+8CC2 <cjk>
	0x48: [`\u8DEF`].string() // U+8DEF <cjk>
	0x49: [`\u9732`].string() // U+9732 <cjk>
	0x4A: [`\u52B4`].string() // U+52B4 <cjk>
	0x4B: [`\u5A41`].string() // U+5A41 <cjk>
	0x4C: [`\u5ECA`].string() // U+5ECA <cjk>
	0x4D: [`\u5F04`].string() // U+5F04 <cjk>
	0x4E: [`\u6717`].string() // U+6717 <cjk>
	0x4F: [`\u697C`].string() // U+697C <cjk>
	0x50: [`\u6994`].string() // U+6994 <cjk>
	0x51: [`\u6D6A`].string() // U+6D6A <cjk>
	0x52: [`\u6F0F`].string() // U+6F0F <cjk>
	0x53: [`\u7262`].string() // U+7262 <cjk>
	0x54: [`\u72FC`].string() // U+72FC <cjk>
	0x55: [`\u7BED`].string() // U+7BED <cjk>
	0x56: [`\u8001`].string() // U+8001 <cjk>
	0x57: [`\u807E`].string() // U+807E <cjk>
	0x58: [`\u874B`].string() // U+874B <cjk>
	0x59: [`\u90CE`].string() // U+90CE <cjk>
	0x5A: [`\u516D`].string() // U+516D <cjk>
	0x5B: [`\u9E93`].string() // U+9E93 <cjk>
	0x5C: [`\u7984`].string() // U+7984 <cjk>
	0x5D: [`\u808B`].string() // U+808B <cjk>
	0x5E: [`\u9332`].string() // U+9332 <cjk>
	0x5F: [`\u8AD6`].string() // U+8AD6 <cjk>
	0x60: [`\u502D`].string() // U+502D <cjk>
	0x61: [`\u548C`].string() // U+548C <cjk>
	0x62: [`\u8A71`].string() // U+8A71 <cjk>
	0x63: [`\u6B6A`].string() // U+6B6A <cjk>
	0x64: [`\u8CC4`].string() // U+8CC4 <cjk>
	0x65: [`\u8107`].string() // U+8107 <cjk>
	0x66: [`\u60D1`].string() // U+60D1 <cjk>
	0x67: [`\u67A0`].string() // U+67A0 <cjk>
	0x68: [`\u9DF2`].string() // U+9DF2 <cjk>
	0x69: [`\u4E99`].string() // U+4E99 <cjk>
	0x6A: [`\u4E98`].string() // U+4E98 <cjk>
	0x6B: [`\u9C10`].string() // U+9C10 <cjk>
	0x6C: [`\u8A6B`].string() // U+8A6B <cjk>
	0x6D: [`\u85C1`].string() // U+85C1 <cjk>
	0x6E: [`\u8568`].string() // U+8568 <cjk>
	0x6F: [`\u6900`].string() // U+6900 <cjk>
	0x70: [`\u6E7E`].string() // U+6E7E <cjk>
	0x71: [`\u7897`].string() // U+7897 <cjk>
	0x72: [`\u8155`].string() // U+8155 <cjk>
	0x73: utf32_to_str(0x20B98) // U+20B9F <cjk>
	0x74: [`\u5B41`].string() // U+5B41 <cjk>
	0x75: [`\u5B56`].string() // U+5B56 <cjk>
	0x76: [`\u5B7D`].string() // U+5B7D <cjk>
	0x77: [`\u5B93`].string() // U+5B93 <cjk>
	0x78: [`\u5BD8`].string() // U+5BD8 <cjk>
	0x79: [`\u5BEC`].string() // U+5BEC <cjk>
	0x7A: [`\u5C12`].string() // U+5C12 <cjk>
	0x7B: [`\u5C1E`].string() // U+5C1E <cjk>
	0x7C: [`\u5C23`].string() // U+5C23 <cjk>
	0x7D: [`\u5C2B`].string() // U+5C2B <cjk>
	0x7E: [`\u378D`].string() // U+378D <cjk>
	0x80: [`\u5C62`].string() // U+5C62 <cjk>
	0x81: [`\uFA3B`].string() // U+FA3B CJK COMPATIBILITY IDEOGRAPH-FA3B
	0x82: [`\uFA3C`].string() // U+FA3C CJK COMPATIBILITY IDEOGRAPH-FA3C
	0x83: utf32_to_str(0x216B4) // U+216B4 <cjk>
	0x84: [`\u5C7A`].string() // U+5C7A <cjk>
	0x85: [`\u5C8F`].string() // U+5C8F <cjk>
	0x86: [`\u5C9F`].string() // U+5C9F <cjk>
	0x87: [`\u5CA3`].string() // U+5CA3 <cjk>
	0x88: [`\u5CAA`].string() // U+5CAA <cjk>
	0x89: [`\u5CBA`].string() // U+5CBA <cjk>
	0x8A: [`\u5CCB`].string() // U+5CCB <cjk>
	0x8B: [`\u5CD0`].string() // U+5CD0 <cjk>
	0x8C: [`\u5CD2`].string() // U+5CD2 <cjk>
	0x8D: [`\u5CF4`].string() // U+5CF4 <cjk>
	0x8E: utf32_to_str(0x21E34) // U+21E34 <cjk>
	0x8F: [`\u37E2`].string() // U+37E2 <cjk>
	0x90: [`\u5D0D`].string() // U+5D0D <cjk>
	0x91: [`\u5D27`].string() // U+5D27 <cjk>
	0x92: [`\uFA11`].string() // U+FA11 CJK COMPATIBILITY IDEOGRAPH-FA11
	0x93: [`\u5D46`].string() // U+5D46 <cjk>
	0x94: [`\u5D47`].string() // U+5D47 <cjk>
	0x95: [`\u5D53`].string() // U+5D53 <cjk>
	0x96: [`\u5D4A`].string() // U+5D4A <cjk>
	0x97: [`\u5D6D`].string() // U+5D6D <cjk>
	0x98: [`\u5D81`].string() // U+5D81 <cjk>
	0x99: [`\u5DA0`].string() // U+5DA0 <cjk>
	0x9A: [`\u5DA4`].string() // U+5DA4 <cjk>
	0x9B: [`\u5DA7`].string() // U+5DA7 <cjk>
	0x9C: [`\u5DB8`].string() // U+5DB8 <cjk>
	0x9D: [`\u5DCB`].string() // U+5DCB <cjk>
	0x9E: [`\u541E`].string() // U+541E <cjk>
	0x9F: [`\u5F0C`].string() // U+5F0C <cjk>
	0xA0: [`\u4E10`].string() // U+4E10 <cjk>
	0xA1: [`\u4E15`].string() // U+4E15 <cjk>
	0xA2: [`\u4E2A`].string() // U+4E2A <cjk>
	0xA3: [`\u4E31`].string() // U+4E31 <cjk>
	0xA4: [`\u4E36`].string() // U+4E36 <cjk>
	0xA5: [`\u4E3C`].string() // U+4E3C <cjk>
	0xA6: [`\u4E3F`].string() // U+4E3F <cjk>
	0xA7: [`\u4E42`].string() // U+4E42 <cjk>
	0xA8: [`\u4E56`].string() // U+4E56 <cjk>
	0xA9: [`\u4E58`].string() // U+4E58 <cjk>
	0xAA: [`\u4E82`].string() // U+4E82 <cjk>
	0xAB: [`\u4E85`].string() // U+4E85 <cjk>
	0xAC: [`\u8C6B`].string() // U+8C6B <cjk>
	0xAD: [`\u4E8A`].string() // U+4E8A <cjk>
	0xAE: [`\u8212`].string() // U+8212 <cjk>
	0xAF: [`\u5F0D`].string() // U+5F0D <cjk>
	0xB0: [`\u4E8E`].string() // U+4E8E <cjk>
	0xB1: [`\u4E9E`].string() // U+4E9E <cjk>
	0xB2: [`\u4E9F`].string() // U+4E9F <cjk>
	0xB3: [`\u4EA0`].string() // U+4EA0 <cjk>
	0xB4: [`\u4EA2`].string() // U+4EA2 <cjk>
	0xB5: [`\u4EB0`].string() // U+4EB0 <cjk>
	0xB6: [`\u4EB3`].string() // U+4EB3 <cjk>
	0xB7: [`\u4EB6`].string() // U+4EB6 <cjk>
	0xB8: [`\u4ECE`].string() // U+4ECE <cjk>
	0xB9: [`\u4ECD`].string() // U+4ECD <cjk>
	0xBA: [`\u4EC4`].string() // U+4EC4 <cjk>
	0xBB: [`\u4EC6`].string() // U+4EC6 <cjk>
	0xBC: [`\u4EC2`].string() // U+4EC2 <cjk>
	0xBD: [`\u4ED7`].string() // U+4ED7 <cjk>
	0xBE: [`\u4EDE`].string() // U+4EDE <cjk>
	0xBF: [`\u4EED`].string() // U+4EED <cjk>
	0xC0: [`\u4EDF`].string() // U+4EDF <cjk>
	0xC1: [`\u4EF7`].string() // U+4EF7 <cjk>
	0xC2: [`\u4F09`].string() // U+4F09 <cjk>
	0xC3: [`\u4F5A`].string() // U+4F5A <cjk>
	0xC4: [`\u4F30`].string() // U+4F30 <cjk>
	0xC5: [`\u4F5B`].string() // U+4F5B <cjk>
	0xC6: [`\u4F5D`].string() // U+4F5D <cjk>
	0xC7: [`\u4F57`].string() // U+4F57 <cjk>
	0xC8: [`\u4F47`].string() // U+4F47 <cjk>
	0xC9: [`\u4F76`].string() // U+4F76 <cjk>
	0xCA: [`\u4F88`].string() // U+4F88 <cjk>
	0xCB: [`\u4F8F`].string() // U+4F8F <cjk>
	0xCC: [`\u4F98`].string() // U+4F98 <cjk>
	0xCD: [`\u4F7B`].string() // U+4F7B <cjk>
	0xCE: [`\u4F69`].string() // U+4F69 <cjk>
	0xCF: [`\u4F70`].string() // U+4F70 <cjk>
	0xD0: [`\u4F91`].string() // U+4F91 <cjk>
	0xD1: [`\u4F6F`].string() // U+4F6F <cjk>
	0xD2: [`\u4F86`].string() // U+4F86 <cjk>
	0xD3: [`\u4F96`].string() // U+4F96 <cjk>
	0xD4: [`\u5118`].string() // U+5118 <cjk>
	0xD5: [`\u4FD4`].string() // U+4FD4 <cjk>
	0xD6: [`\u4FDF`].string() // U+4FDF <cjk>
	0xD7: [`\u4FCE`].string() // U+4FCE <cjk>
	0xD8: [`\u4FD8`].string() // U+4FD8 <cjk>
	0xD9: [`\u4FDB`].string() // U+4FDB <cjk>
	0xDA: [`\u4FD1`].string() // U+4FD1 <cjk>
	0xDB: [`\u4FDA`].string() // U+4FDA <cjk>
	0xDC: [`\u4FD0`].string() // U+4FD0 <cjk>
	0xDD: [`\u4FE4`].string() // U+4FE4 <cjk>
	0xDE: [`\u4FE5`].string() // U+4FE5 <cjk>
	0xDF: [`\u501A`].string() // U+501A <cjk>
	0xE0: [`\u5028`].string() // U+5028 <cjk>
	0xE1: [`\u5014`].string() // U+5014 <cjk>
	0xE2: [`\u502A`].string() // U+502A <cjk>
	0xE3: [`\u5025`].string() // U+5025 <cjk>
	0xE4: [`\u5005`].string() // U+5005 <cjk>
	0xE5: [`\u4F1C`].string() // U+4F1C <cjk>
	0xE6: [`\u4FF6`].string() // U+4FF6 <cjk>
	0xE7: [`\u5021`].string() // U+5021 <cjk>
	0xE8: [`\u5029`].string() // U+5029 <cjk>
	0xE9: [`\u502C`].string() // U+502C <cjk>
	0xEA: [`\u4FFE`].string() // U+4FFE <cjk>
	0xEB: [`\u4FEF`].string() // U+4FEF <cjk>
	0xEC: [`\u5011`].string() // U+5011 <cjk>
	0xED: [`\u5006`].string() // U+5006 <cjk>
	0xEE: [`\u5043`].string() // U+5043 <cjk>
	0xEF: [`\u5047`].string() // U+5047 <cjk>
	0xF0: [`\u6703`].string() // U+6703 <cjk>
	0xF1: [`\u5055`].string() // U+5055 <cjk>
	0xF2: [`\u5050`].string() // U+5050 <cjk>
	0xF3: [`\u5048`].string() // U+5048 <cjk>
	0xF4: [`\u505A`].string() // U+505A <cjk>
	0xF5: [`\u5056`].string() // U+5056 <cjk>
	0xF6: [`\u506C`].string() // U+506C <cjk>
	0xF7: [`\u5078`].string() // U+5078 <cjk>
	0xF8: [`\u5080`].string() // U+5080 <cjk>
	0xF9: [`\u509A`].string() // U+509A <cjk>
	0xFA: [`\u5085`].string() // U+5085 <cjk>
	0xFB: [`\u50B4`].string() // U+50B4 <cjk>
	0xFC: [`\u50B2`].string() // U+50B2 <cjk>
}

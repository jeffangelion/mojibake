module mojibake

const jis_x_0213_doublebyte_0x86 = {
	0x40: [`\u0294`].string() // U+0294 LATIN LETTER GLOTTAL STOP
	0x41: [`\u0266`].string() // U+0266 LATIN SMALL LETTER H WITH HOOK
	0x42: [`\u0298`].string() // U+0298 LATIN LETTER BILABIAL CLICK
	0x43: [`\u01C2`].string() // U+01C2 LATIN LETTER ALVEOLAR CLICK
	0x44: [`\u0253`].string() // U+0253 LATIN SMALL LETTER B WITH HOOK
	0x45: [`\u0257`].string() // U+0257 LATIN SMALL LETTER D WITH HOOK
	0x46: [`\u0284`].string() // U+0284 LATIN SMALL LETTER DOTLESS J WITH STROKE AND HOOK
	0x47: [`\u0260`].string() // U+0260 LATIN SMALL LETTER G WITH HOOK
	0x48: [`\u0193`].string() // U+0193 LATIN CAPITAL LETTER G WITH HOOK
	0x49: [`\u0153`].string() // U+0153 LATIN SMALL LIGATURE OE
	0x4A: [`\u0152`].string() // U+0152 LATIN CAPITAL LIGATURE OE
	0x4B: [`\u0268`].string() // U+0268 LATIN SMALL LETTER I WITH STROKE
	0x4C: [`\u0289`].string() // U+0289 LATIN SMALL LETTER U BAR
	0x4D: [`\u0258`].string() // U+0258 LATIN SMALL LETTER REVERSED E
	0x4E: [`\u0275`].string() // U+0275 LATIN SMALL LETTER BARRED O
	0x4F: [`\u0259`].string() // U+0259 LATIN SMALL LETTER SCHWA
	0x50: [`\u025C`].string() // U+025C LATIN SMALL LETTER REVERSED OPEN E
	0x51: [`\u025E`].string() // U+025E LATIN SMALL LETTER CLOSED REVERSED OPEN E
	0x52: [`\u0250`].string() // U+0250 LATIN SMALL LETTER TURNED A
	0x53: [`\u026F`].string() // U+026F LATIN SMALL LETTER TURNED M
	0x54: [`\u028A`].string() // U+028A LATIN SMALL LETTER UPSILON
	0x55: [`\u0264`].string() // U+0264 LATIN SMALL LETTER RAMS HORN
	0x56: [`\u028C`].string() // U+028C LATIN SMALL LETTER TURNED V
	0x57: [`\u0254`].string() // U+0254 LATIN SMALL LETTER OPEN O
	0x58: [`\u0251`].string() // U+0251 LATIN SMALL LETTER ALPHA
	0x59: [`\u0252`].string() // U+0252 LATIN SMALL LETTER TURNED ALPHA
	0x5A: [`\u028D`].string() // U+028D LATIN SMALL LETTER TURNED W
	0x5B: [`\u0265`].string() // U+0265 LATIN SMALL LETTER TURNED H
	0x5C: [`\u02A2`].string() // U+02A2 LATIN LETTER REVERSED GLOTTAL STOP WITH STROKE
	0x5D: [`\u02A1`].string() // U+02A1 LATIN LETTER GLOTTAL STOP WITH STROKE
	0x5E: [`\u0255`].string() // U+0255 LATIN SMALL LETTER C WITH CURL
	0x5F: [`\u0291`].string() // U+0291 LATIN SMALL LETTER Z WITH CURL
	0x60: [`\u027A`].string() // U+027A LATIN SMALL LETTER TURNED R WITH LONG LEG
	0x61: [`\u0267`].string() // U+0267 LATIN SMALL LETTER HENG WITH HOOK
	0x62: [`\u025A`].string() // U+025A LATIN SMALL LETTER SCHWA WITH HOOK
	0x63: [`\u00E6`,`\u0300`].string() // U+00E6+0300
	0x64: [`\u01FD`].string() // U+01FD LATIN SMALL LETTER AE WITH ACUTE
	0x65: [`\u1F70`].string() // U+1F70 GREEK SMALL LETTER ALPHA WITH VARIA
	0x66: [`\u1F71`].string() // U+1F71 GREEK SMALL LETTER ALPHA WITH OXIA
	0x67: [`\u0254`,`\u0300`].string() // U+0254+0300
	0x68: [`\u0254`,`\u0301`].string() // U+0254+0301
	0x69: [`\u028C`,`\u0300`].string() // U+028C+0300
	0x6A: [`\u028C`,`\u0301`].string() // U+028C+0301
	0x6B: [`\u0259`,`\u0300`].string() // U+0259+0300
	0x6C: [`\u0259`,`\u0301`].string() // U+0259+0301
	0x6D: [`\u025A`,`\u0300`].string() // U+025A+0300
	0x6E: [`\u025A`,`\u0301`].string() // U+025A+0301
	0x6F: [`\u1F72`].string() // U+1F72 GREEK SMALL LETTER EPSILON WITH VARIA
	0x70: [`\u1F73`].string() // U+1F73 GREEK SMALL LETTER EPSILON WITH OXIA
	0x71: [`\u0361`].string() // U+0361 COMBINING DOUBLE INVERTED BREVE
	0x72: [`\u02C8`].string() // U+02C8 MODIFIER LETTER VERTICAL LINE
	0x73: [`\u02CC`].string() // U+02CC MODIFIER LETTER LOW VERTICAL LINE
	0x74: [`\u02D0`].string() // U+02D0 MODIFIER LETTER TRIANGULAR COLON
	0x75: [`\u02D1`].string() // U+02D1 MODIFIER LETTER HALF TRIANGULAR COLON
	0x76: [`\u0306`].string() // U+0306 COMBINING BREVE
	0x77: [`\u203F`].string() // U+203F UNDERTIE
	0x78: [`\u030B`].string() // U+030B COMBINING DOUBLE ACUTE ACCENT
	0x79: [`\u0301`].string() // U+0301 COMBINING ACUTE ACCENT
	0x7A: [`\u0304`].string() // U+0304 COMBINING MACRON
	0x7B: [`\u0300`].string() // U+0300 COMBINING GRAVE ACCENT
	0x7C: [`\u030F`].string() // U+030F COMBINING DOUBLE GRAVE ACCENT
	0x7D: [`\u030C`].string() // U+030C COMBINING CARON
	0x7E: [`\u0302`].string() // U+0302 COMBINING CIRCUMFLEX ACCENT
	0x80: [`\u02E5`].string() // U+02E5 MODIFIER LETTER EXTRA-HIGH TONE BAR
	0x81: [`\u02E6`].string() // U+02E6 MODIFIER LETTER HIGH TONE BAR
	0x82: [`\u02E7`].string() // U+02E7 MODIFIER LETTER MID TONE BAR
	0x83: [`\u02E8`].string() // U+02E8 MODIFIER LETTER LOW TONE BAR
	0x84: [`\u02E9`].string() // U+02E9 MODIFIER LETTER EXTRA-LOW TONE BAR
	0x85: [`\u02E9`,`\u02E5`].string() // U+02E9+02E5
	0x86: [`\u02E5`,`\u02E9`].string() // U+02E5+02E9
	0x87: [`\u0325`].string() // U+0325 COMBINING RING BELOW
	0x88: [`\u032C`].string() // U+032C COMBINING CARON BELOW
	0x89: [`\u0339`].string() // U+0339 COMBINING RIGHT HALF RING BELOW
	0x8A: [`\u031C`].string() // U+031C COMBINING LEFT HALF RING BELOW
	0x8B: [`\u031F`].string() // U+031F COMBINING PLUS SIGN BELOW
	0x8C: [`\u0320`].string() // U+0320 COMBINING MINUS SIGN BELOW
	0x8D: [`\u0308`].string() // U+0308 COMBINING DIAERESIS
	0x8E: [`\u033D`].string() // U+033D COMBINING X ABOVE
	0x8F: [`\u0329`].string() // U+0329 COMBINING VERTICAL LINE BELOW
	0x90: [`\u032F`].string() // U+032F COMBINING INVERTED BREVE BELOW
	0x91: [`\u02DE`].string() // U+02DE MODIFIER LETTER RHOTIC HOOK
	0x92: [`\u0324`].string() // U+0324 COMBINING DIAERESIS BELOW
	0x93: [`\u0330`].string() // U+0330 COMBINING TILDE BELOW
	0x94: [`\u033C`].string() // U+033C COMBINING SEAGULL BELOW
	0x95: [`\u0334`].string() // U+0334 COMBINING TILDE OVERLAY
	0x96: [`\u031D`].string() // U+031D COMBINING UP TACK BELOW
	0x97: [`\u031E`].string() // U+031E COMBINING DOWN TACK BELOW
	0x98: [`\u0318`].string() // U+0318 COMBINING LEFT TACK BELOW
	0x99: [`\u0319`].string() // U+0319 COMBINING RIGHT TACK BELOW
	0x9A: [`\u032A`].string() // U+032A COMBINING BRIDGE BELOW
	0x9B: [`\u033A`].string() // U+033A COMBINING INVERTED BRIDGE BELOW
	0x9C: [`\u033B`].string() // U+033B COMBINING SQUARE BELOW
	0x9D: [`\u0303`].string() // U+0303 COMBINING TILDE
	0x9E: [`\u031A`].string() // U+031A COMBINING LEFT ANGLE ABOVE
	0x9F: [`\u2776`].string() // U+2776 DINGBAT NEGATIVE CIRCLED DIGIT ONE
	0xA0: [`\u2777`].string() // U+2777 DINGBAT NEGATIVE CIRCLED DIGIT TWO
	0xA1: [`\u2778`].string() // U+2778 DINGBAT NEGATIVE CIRCLED DIGIT THREE
	0xA2: [`\u2779`].string() // U+2779 DINGBAT NEGATIVE CIRCLED DIGIT FOUR
	0xA3: [`\u277A`].string() // U+277A DINGBAT NEGATIVE CIRCLED DIGIT FIVE
	0xA4: [`\u277B`].string() // U+277B DINGBAT NEGATIVE CIRCLED DIGIT SIX
	0xA5: [`\u277C`].string() // U+277C DINGBAT NEGATIVE CIRCLED DIGIT SEVEN
	0xA6: [`\u277D`].string() // U+277D DINGBAT NEGATIVE CIRCLED DIGIT EIGHT
	0xA7: [`\u277E`].string() // U+277E DINGBAT NEGATIVE CIRCLED DIGIT NINE
	0xA8: [`\u277F`].string() // U+277F DINGBAT NEGATIVE CIRCLED NUMBER TEN
	0xA9: [`\u24EB`].string() // U+24EB NEGATIVE CIRCLED NUMBER ELEVEN
	0xAA: [`\u24EC`].string() // U+24EC NEGATIVE CIRCLED NUMBER TWELVE
	0xAB: [`\u24ED`].string() // U+24ED NEGATIVE CIRCLED NUMBER THIRTEEN
	0xAC: [`\u24EE`].string() // U+24EE NEGATIVE CIRCLED NUMBER FOURTEEN
	0xAD: [`\u24EF`].string() // U+24EF NEGATIVE CIRCLED NUMBER FIFTEEN
	0xAE: [`\u24F0`].string() // U+24F0 NEGATIVE CIRCLED NUMBER SIXTEEN
	0xAF: [`\u24F1`].string() // U+24F1 NEGATIVE CIRCLED NUMBER SEVENTEEN
	0xB0: [`\u24F2`].string() // U+24F2 NEGATIVE CIRCLED NUMBER EIGHTEEN
	0xB1: [`\u24F3`].string() // U+24F3 NEGATIVE CIRCLED NUMBER NINETEEN
	0xB2: [`\u24F4`].string() // U+24F4 NEGATIVE CIRCLED NUMBER TWENTY
	0xB3: [`\u2170`].string() // U+2170 SMALL ROMAN NUMERAL ONE
	0xB4: [`\u2171`].string() // U+2171 SMALL ROMAN NUMERAL TWO
	0xB5: [`\u2172`].string() // U+2172 SMALL ROMAN NUMERAL THREE
	0xB6: [`\u2173`].string() // U+2173 SMALL ROMAN NUMERAL FOUR
	0xB7: [`\u2174`].string() // U+2174 SMALL ROMAN NUMERAL FIVE
	0xB8: [`\u2175`].string() // U+2175 SMALL ROMAN NUMERAL SIX
	0xB9: [`\u2176`].string() // U+2176 SMALL ROMAN NUMERAL SEVEN
	0xBA: [`\u2177`].string() // U+2177 SMALL ROMAN NUMERAL EIGHT
	0xBB: [`\u2178`].string() // U+2178 SMALL ROMAN NUMERAL NINE
	0xBC: [`\u2179`].string() // U+2179 SMALL ROMAN NUMERAL TEN
	0xBD: [`\u217A`].string() // U+217A SMALL ROMAN NUMERAL ELEVEN
	0xBE: [`\u217B`].string() // U+217B SMALL ROMAN NUMERAL TWELVE
	0xBF: [`\u24D0`].string() // U+24D0 CIRCLED LATIN SMALL LETTER A
	0xC0: [`\u24D1`].string() // U+24D1 CIRCLED LATIN SMALL LETTER B
	0xC1: [`\u24D2`].string() // U+24D2 CIRCLED LATIN SMALL LETTER C
	0xC2: [`\u24D3`].string() // U+24D3 CIRCLED LATIN SMALL LETTER D
	0xC3: [`\u24D4`].string() // U+24D4 CIRCLED LATIN SMALL LETTER E
	0xC4: [`\u24D5`].string() // U+24D5 CIRCLED LATIN SMALL LETTER F
	0xC5: [`\u24D6`].string() // U+24D6 CIRCLED LATIN SMALL LETTER G
	0xC6: [`\u24D7`].string() // U+24D7 CIRCLED LATIN SMALL LETTER H
	0xC7: [`\u24D8`].string() // U+24D8 CIRCLED LATIN SMALL LETTER I
	0xC8: [`\u24D9`].string() // U+24D9 CIRCLED LATIN SMALL LETTER J
	0xC9: [`\u24DA`].string() // U+24DA CIRCLED LATIN SMALL LETTER K
	0xCA: [`\u24DB`].string() // U+24DB CIRCLED LATIN SMALL LETTER L
	0xCB: [`\u24DC`].string() // U+24DC CIRCLED LATIN SMALL LETTER M
	0xCC: [`\u24DD`].string() // U+24DD CIRCLED LATIN SMALL LETTER N
	0xCD: [`\u24DE`].string() // U+24DE CIRCLED LATIN SMALL LETTER O
	0xCE: [`\u24DF`].string() // U+24DF CIRCLED LATIN SMALL LETTER P
	0xCF: [`\u24E0`].string() // U+24E0 CIRCLED LATIN SMALL LETTER Q
	0xD0: [`\u24E1`].string() // U+24E1 CIRCLED LATIN SMALL LETTER R
	0xD1: [`\u24E2`].string() // U+24E2 CIRCLED LATIN SMALL LETTER S
	0xD2: [`\u24E3`].string() // U+24E3 CIRCLED LATIN SMALL LETTER T
	0xD3: [`\u24E4`].string() // U+24E4 CIRCLED LATIN SMALL LETTER U
	0xD4: [`\u24E5`].string() // U+24E5 CIRCLED LATIN SMALL LETTER V
	0xD5: [`\u24E6`].string() // U+24E6 CIRCLED LATIN SMALL LETTER W
	0xD6: [`\u24E7`].string() // U+24E7 CIRCLED LATIN SMALL LETTER X
	0xD7: [`\u24E8`].string() // U+24E8 CIRCLED LATIN SMALL LETTER Y
	0xD8: [`\u24E9`].string() // U+24E9 CIRCLED LATIN SMALL LETTER Z
	0xD9: [`\u32D0`].string() // U+32D0 CIRCLED KATAKANA A
	0xDA: [`\u32D1`].string() // U+32D1 CIRCLED KATAKANA I
	0xDB: [`\u32D2`].string() // U+32D2 CIRCLED KATAKANA U
	0xDC: [`\u32D3`].string() // U+32D3 CIRCLED KATAKANA E
	0xDD: [`\u32D4`].string() // U+32D4 CIRCLED KATAKANA O
	0xDE: [`\u32D5`].string() // U+32D5 CIRCLED KATAKANA KA
	0xDF: [`\u32D6`].string() // U+32D6 CIRCLED KATAKANA KI
	0xE0: [`\u32D7`].string() // U+32D7 CIRCLED KATAKANA KU
	0xE1: [`\u32D8`].string() // U+32D8 CIRCLED KATAKANA KE
	0xE2: [`\u32D9`].string() // U+32D9 CIRCLED KATAKANA KO
	0xE3: [`\u32DA`].string() // U+32DA CIRCLED KATAKANA SA
	0xE4: [`\u32DB`].string() // U+32DB CIRCLED KATAKANA SI
	0xE5: [`\u32DC`].string() // U+32DC CIRCLED KATAKANA SU
	0xE6: [`\u32DD`].string() // U+32DD CIRCLED KATAKANA SE
	0xE7: [`\u32DE`].string() // U+32DE CIRCLED KATAKANA SO
	0xE8: [`\u32DF`].string() // U+32DF CIRCLED KATAKANA TA
	0xE9: [`\u32E0`].string() // U+32E0 CIRCLED KATAKANA TI
	0xEA: [`\u32E1`].string() // U+32E1 CIRCLED KATAKANA TU
	0xEB: [`\u32E2`].string() // U+32E2 CIRCLED KATAKANA TE
	0xEC: [`\u32E3`].string() // U+32E3 CIRCLED KATAKANA TO
	0xED: [`\u32FA`].string() // U+32FA CIRCLED KATAKANA RO
	0xEE: [`\u32E9`].string() // U+32E9 CIRCLED KATAKANA HA
	0xEF: [`\u32E5`].string() // U+32E5 CIRCLED KATAKANA NI
	0xF0: [`\u32ED`].string() // U+32ED CIRCLED KATAKANA HO
	0xF1: [`\u32EC`].string() // U+32EC CIRCLED KATAKANA HE
	0xFB: [`\u2051`].string() // U+2051 TWO ASTERISKS ALIGNED VERTICALLY
	0xFC: [`\u2042`].string() // U+2042 ASTERISM
}

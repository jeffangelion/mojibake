module mojibake

const jis_x_0213_doublebyte_0x96 = {
	0x40: [`\u6CD5`].string() // U+6CD5 <cjk>
	0x41: [`\u6CE1`].string() // U+6CE1 <cjk>
	0x42: [`\u70F9`].string() // U+70F9 <cjk>
	0x43: [`\u7832`].string() // U+7832 <cjk>
	0x44: [`\u7E2B`].string() // U+7E2B <cjk>
	0x45: [`\u80DE`].string() // U+80DE <cjk>
	0x46: [`\u82B3`].string() // U+82B3 <cjk>
	0x47: [`\u840C`].string() // U+840C <cjk>
	0x48: [`\u84EC`].string() // U+84EC <cjk>
	0x49: [`\u8702`].string() // U+8702 <cjk>
	0x4A: [`\u8912`].string() // U+8912 <cjk>
	0x4B: [`\u8A2A`].string() // U+8A2A <cjk>
	0x4C: [`\u8C4A`].string() // U+8C4A <cjk>
	0x4D: [`\u90A6`].string() // U+90A6 <cjk>
	0x4E: [`\u92D2`].string() // U+92D2 <cjk>
	0x4F: [`\u98FD`].string() // U+98FD <cjk>
	0x50: [`\u9CF3`].string() // U+9CF3 <cjk>
	0x51: [`\u9D6C`].string() // U+9D6C <cjk>
	0x52: [`\u4E4F`].string() // U+4E4F <cjk>
	0x53: [`\u4EA1`].string() // U+4EA1 <cjk>
	0x54: [`\u508D`].string() // U+508D <cjk>
	0x55: [`\u5256`].string() // U+5256 <cjk>
	0x56: [`\u574A`].string() // U+574A <cjk>
	0x57: [`\u59A8`].string() // U+59A8 <cjk>
	0x58: [`\u5E3D`].string() // U+5E3D <cjk>
	0x59: [`\u5FD8`].string() // U+5FD8 <cjk>
	0x5A: [`\u5FD9`].string() // U+5FD9 <cjk>
	0x5B: [`\u623F`].string() // U+623F <cjk>
	0x5C: [`\u66B4`].string() // U+66B4 <cjk>
	0x5D: [`\u671B`].string() // U+671B <cjk>
	0x5E: [`\u67D0`].string() // U+67D0 <cjk>
	0x5F: [`\u68D2`].string() // U+68D2 <cjk>
	0x60: [`\u5192`].string() // U+5192 <cjk>
	0x61: [`\u7D21`].string() // U+7D21 <cjk>
	0x62: [`\u80AA`].string() // U+80AA <cjk>
	0x63: [`\u81A8`].string() // U+81A8 <cjk>
	0x64: [`\u8B00`].string() // U+8B00 <cjk>
	0x65: [`\u8C8C`].string() // U+8C8C <cjk>
	0x66: [`\u8CBF`].string() // U+8CBF <cjk>
	0x67: [`\u927E`].string() // U+927E <cjk>
	0x68: [`\u9632`].string() // U+9632 <cjk>
	0x69: [`\u5420`].string() // U+5420 <cjk>
	0x6A: [`\u982C`].string() // U+982C <cjk>
	0x6B: [`\u5317`].string() // U+5317 <cjk>
	0x6C: [`\u50D5`].string() // U+50D5 <cjk>
	0x6D: [`\u535C`].string() // U+535C <cjk>
	0x6E: [`\u58A8`].string() // U+58A8 <cjk>
	0x6F: [`\u64B2`].string() // U+64B2 <cjk>
	0x70: [`\u6734`].string() // U+6734 <cjk>
	0x71: [`\u7267`].string() // U+7267 <cjk>
	0x72: [`\u7766`].string() // U+7766 <cjk>
	0x73: [`\u7A46`].string() // U+7A46 <cjk>
	0x74: [`\u91E6`].string() // U+91E6 <cjk>
	0x75: [`\u52C3`].string() // U+52C3 <cjk>
	0x76: [`\u6CA1`].string() // U+6CA1 <cjk>
	0x77: [`\u6B86`].string() // U+6B86 <cjk>
	0x78: [`\u5800`].string() // U+5800 <cjk>
	0x79: [`\u5E4C`].string() // U+5E4C <cjk>
	0x7A: [`\u5954`].string() // U+5954 <cjk>
	0x7B: [`\u672C`].string() // U+672C <cjk>
	0x7C: [`\u7FFB`].string() // U+7FFB <cjk>
	0x7D: [`\u51E1`].string() // U+51E1 <cjk>
	0x7E: [`\u76C6`].string() // U+76C6 <cjk>
	0x80: [`\u6469`].string() // U+6469 <cjk>
	0x81: [`\u78E8`].string() // U+78E8 <cjk>
	0x82: [`\u9B54`].string() // U+9B54 <cjk>
	0x83: [`\u9EBB`].string() // U+9EBB <cjk>
	0x84: [`\u57CB`].string() // U+57CB <cjk>
	0x85: [`\u59B9`].string() // U+59B9 <cjk>
	0x86: [`\u6627`].string() // U+6627 <cjk>
	0x87: [`\u679A`].string() // U+679A <cjk>
	0x88: [`\u6BCE`].string() // U+6BCE <cjk>
	0x89: [`\u54E9`].string() // U+54E9 <cjk>
	0x8A: [`\u69D9`].string() // U+69D9 <cjk>
	0x8B: [`\u5E55`].string() // U+5E55 <cjk>
	0x8C: [`\u819C`].string() // U+819C <cjk>
	0x8D: [`\u6795`].string() // U+6795 <cjk>
	0x8E: [`\u9BAA`].string() // U+9BAA <cjk>
	0x8F: [`\u67FE`].string() // U+67FE <cjk>
	0x90: [`\u9C52`].string() // U+9C52 <cjk>
	0x91: [`\u685D`].string() // U+685D <cjk>
	0x92: [`\u4EA6`].string() // U+4EA6 <cjk>
	0x93: [`\u4FE3`].string() // U+4FE3 <cjk>
	0x94: [`\u53C8`].string() // U+53C8 <cjk>
	0x95: [`\u62B9`].string() // U+62B9 <cjk>
	0x96: [`\u672B`].string() // U+672B <cjk>
	0x97: [`\u6CAB`].string() // U+6CAB <cjk>
	0x98: [`\u8FC4`].string() // U+8FC4 <cjk>
	0x99: [`\u4FAD`].string() // U+4FAD <cjk>
	0x9A: [`\u7E6D`].string() // U+7E6D <cjk>
	0x9B: [`\u9EBF`].string() // U+9EBF <cjk>
	0x9C: [`\u4E07`].string() // U+4E07 <cjk>
	0x9D: [`\u6162`].string() // U+6162 <cjk>
	0x9E: [`\u6E80`].string() // U+6E80 <cjk>
	0x9F: [`\u6F2B`].string() // U+6F2B <cjk>
	0xA0: [`\u8513`].string() // U+8513 <cjk>
	0xA1: [`\u5473`].string() // U+5473 <cjk>
	0xA2: [`\u672A`].string() // U+672A <cjk>
	0xA3: [`\u9B45`].string() // U+9B45 <cjk>
	0xA4: [`\u5DF3`].string() // U+5DF3 <cjk>
	0xA5: [`\u7B95`].string() // U+7B95 <cjk>
	0xA6: [`\u5CAC`].string() // U+5CAC <cjk>
	0xA7: [`\u5BC6`].string() // U+5BC6 <cjk>
	0xA8: [`\u871C`].string() // U+871C <cjk>
	0xA9: [`\u6E4A`].string() // U+6E4A <cjk>
	0xAA: [`\u84D1`].string() // U+84D1 <cjk>
	0xAB: [`\u7A14`].string() // U+7A14 <cjk>
	0xAC: [`\u8108`].string() // U+8108 <cjk>
	0xAD: [`\u5999`].string() // U+5999 <cjk>
	0xAE: [`\u7C8D`].string() // U+7C8D <cjk>
	0xAF: [`\u6C11`].string() // U+6C11 <cjk>
	0xB0: [`\u7720`].string() // U+7720 <cjk>
	0xB1: [`\u52D9`].string() // U+52D9 <cjk>
	0xB2: [`\u5922`].string() // U+5922 <cjk>
	0xB3: [`\u7121`].string() // U+7121 <cjk>
	0xB4: [`\u725F`].string() // U+725F <cjk>
	0xB5: [`\u77DB`].string() // U+77DB <cjk>
	0xB6: [`\u9727`].string() // U+9727 <cjk>
	0xB7: [`\u9D61`].string() // U+9D61 <cjk>
	0xB8: [`\u690B`].string() // U+690B <cjk>
	0xB9: [`\u5A7F`].string() // U+5A7F <cjk>
	0xBA: [`\u5A18`].string() // U+5A18 <cjk>
	0xBB: [`\u51A5`].string() // U+51A5 <cjk>
	0xBC: [`\u540D`].string() // U+540D <cjk>
	0xBD: [`\u547D`].string() // U+547D <cjk>
	0xBE: [`\u660E`].string() // U+660E <cjk>
	0xBF: [`\u76DF`].string() // U+76DF <cjk>
	0xC0: [`\u8FF7`].string() // U+8FF7 <cjk>
	0xC1: [`\u9298`].string() // U+9298 <cjk>
	0xC2: [`\u9CF4`].string() // U+9CF4 <cjk>
	0xC3: [`\u59EA`].string() // U+59EA <cjk>
	0xC4: [`\u725D`].string() // U+725D <cjk>
	0xC5: [`\u6EC5`].string() // U+6EC5 <cjk>
	0xC6: [`\u514D`].string() // U+514D <cjk>
	0xC7: [`\u68C9`].string() // U+68C9 <cjk>
	0xC8: [`\u7DBF`].string() // U+7DBF <cjk>
	0xC9: [`\u7DEC`].string() // U+7DEC <cjk>
	0xCA: [`\u9762`].string() // U+9762 <cjk>
	0xCB: [`\u9EBA`].string() // U+9EBA <cjk>
	0xCC: [`\u6478`].string() // U+6478 <cjk>
	0xCD: [`\u6A21`].string() // U+6A21 <cjk>
	0xCE: [`\u8302`].string() // U+8302 <cjk>
	0xCF: [`\u5984`].string() // U+5984 <cjk>
	0xD0: [`\u5B5F`].string() // U+5B5F <cjk>
	0xD1: [`\u6BDB`].string() // U+6BDB <cjk>
	0xD2: [`\u731B`].string() // U+731B <cjk>
	0xD3: [`\u76F2`].string() // U+76F2 <cjk>
	0xD4: [`\u7DB2`].string() // U+7DB2 <cjk>
	0xD5: [`\u8017`].string() // U+8017 <cjk>
	0xD6: [`\u8499`].string() // U+8499 <cjk>
	0xD7: [`\u5132`].string() // U+5132 <cjk>
	0xD8: [`\u6728`].string() // U+6728 <cjk>
	0xD9: [`\u9ED9`].string() // U+9ED9 <cjk>
	0xDA: [`\u76EE`].string() // U+76EE <cjk>
	0xDB: [`\u6762`].string() // U+6762 <cjk>
	0xDC: [`\u52FF`].string() // U+52FF <cjk>
	0xDD: [`\u9905`].string() // U+9905 <cjk>
	0xDE: [`\u5C24`].string() // U+5C24 <cjk>
	0xDF: [`\u623B`].string() // U+623B <cjk>
	0xE0: [`\u7C7E`].string() // U+7C7E <cjk>
	0xE1: [`\u8CB0`].string() // U+8CB0 <cjk>
	0xE2: [`\u554F`].string() // U+554F <cjk>
	0xE3: [`\u60B6`].string() // U+60B6 <cjk>
	0xE4: [`\u7D0B`].string() // U+7D0B <cjk>
	0xE5: [`\u9580`].string() // U+9580 <cjk>
	0xE6: [`\u5301`].string() // U+5301 <cjk>
	0xE7: [`\u4E5F`].string() // U+4E5F <cjk>
	0xE8: [`\u51B6`].string() // U+51B6 <cjk>
	0xE9: [`\u591C`].string() // U+591C <cjk>
	0xEA: [`\u723A`].string() // U+723A <cjk>
	0xEB: [`\u8036`].string() // U+8036 <cjk>
	0xEC: [`\u91CE`].string() // U+91CE <cjk>
	0xED: [`\u5F25`].string() // U+5F25 <cjk>
	0xEE: [`\u77E2`].string() // U+77E2 <cjk>
	0xEF: [`\u5384`].string() // U+5384 <cjk>
	0xF0: [`\u5F79`].string() // U+5F79 <cjk>
	0xF1: [`\u7D04`].string() // U+7D04 <cjk>
	0xF2: [`\u85AC`].string() // U+85AC <cjk>
	0xF3: [`\u8A33`].string() // U+8A33 <cjk>
	0xF4: [`\u8E8D`].string() // U+8E8D <cjk>
	0xF5: [`\u9756`].string() // U+9756 <cjk>
	0xF6: [`\u67F3`].string() // U+67F3 <cjk>
	0xF7: [`\u85AE`].string() // U+85AE <cjk>
	0xF8: [`\u9453`].string() // U+9453 <cjk>
	0xF9: [`\u6109`].string() // U+6109 <cjk>
	0xFA: [`\u6108`].string() // U+6108 <cjk>
	0xFB: [`\u6CB9`].string() // U+6CB9 <cjk>
	0xFC: [`\u7652`].string() // U+7652 <cjk>
}

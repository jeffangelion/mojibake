module mojibake

const jis_x_0213_doublebyte_0x8d = {
	0x40: [`\u540E`].string() // U+540E <cjk>
	0x41: [`\u5589`].string() // U+5589 <cjk>
	0x42: [`\u5751`].string() // U+5751 <cjk>
	0x43: [`\u57A2`].string() // U+57A2 <cjk>
	0x44: [`\u597D`].string() // U+597D <cjk>
	0x45: [`\u5B54`].string() // U+5B54 <cjk>
	0x46: [`\u5B5D`].string() // U+5B5D <cjk>
	0x47: [`\u5B8F`].string() // U+5B8F <cjk>
	0x48: [`\u5DE5`].string() // U+5DE5 <cjk>
	0x49: [`\u5DE7`].string() // U+5DE7 <cjk>
	0x4A: [`\u5DF7`].string() // U+5DF7 <cjk>
	0x4B: [`\u5E78`].string() // U+5E78 <cjk>
	0x4C: [`\u5E83`].string() // U+5E83 <cjk>
	0x4D: [`\u5E9A`].string() // U+5E9A <cjk>
	0x4E: [`\u5EB7`].string() // U+5EB7 <cjk>
	0x4F: [`\u5F18`].string() // U+5F18 <cjk>
	0x50: [`\u6052`].string() // U+6052 <cjk>
	0x51: [`\u614C`].string() // U+614C <cjk>
	0x52: [`\u6297`].string() // U+6297 <cjk>
	0x53: [`\u62D8`].string() // U+62D8 <cjk>
	0x54: [`\u63A7`].string() // U+63A7 <cjk>
	0x55: [`\u653B`].string() // U+653B <cjk>
	0x56: [`\u6602`].string() // U+6602 <cjk>
	0x57: [`\u6643`].string() // U+6643 <cjk>
	0x58: [`\u66F4`].string() // U+66F4 <cjk>
	0x59: [`\u676D`].string() // U+676D <cjk>
	0x5A: [`\u6821`].string() // U+6821 <cjk>
	0x5B: [`\u6897`].string() // U+6897 <cjk>
	0x5C: [`\u69CB`].string() // U+69CB <cjk>
	0x5D: [`\u6C5F`].string() // U+6C5F <cjk>
	0x5E: [`\u6D2A`].string() // U+6D2A <cjk>
	0x5F: [`\u6D69`].string() // U+6D69 <cjk>
	0x60: [`\u6E2F`].string() // U+6E2F <cjk>
	0x61: [`\u6E9D`].string() // U+6E9D <cjk>
	0x62: [`\u7532`].string() // U+7532 <cjk>
	0x63: [`\u7687`].string() // U+7687 <cjk>
	0x64: [`\u786C`].string() // U+786C <cjk>
	0x65: [`\u7A3F`].string() // U+7A3F <cjk>
	0x66: [`\u7CE0`].string() // U+7CE0 <cjk>
	0x67: [`\u7D05`].string() // U+7D05 <cjk>
	0x68: [`\u7D18`].string() // U+7D18 <cjk>
	0x69: [`\u7D5E`].string() // U+7D5E <cjk>
	0x6A: [`\u7DB1`].string() // U+7DB1 <cjk>
	0x6B: [`\u8015`].string() // U+8015 <cjk>
	0x6C: [`\u8003`].string() // U+8003 <cjk>
	0x6D: [`\u80AF`].string() // U+80AF <cjk>
	0x6E: [`\u80B1`].string() // U+80B1 <cjk>
	0x6F: [`\u8154`].string() // U+8154 <cjk>
	0x70: [`\u818F`].string() // U+818F <cjk>
	0x71: [`\u822A`].string() // U+822A <cjk>
	0x72: [`\u8352`].string() // U+8352 <cjk>
	0x73: [`\u884C`].string() // U+884C <cjk>
	0x74: [`\u8861`].string() // U+8861 <cjk>
	0x75: [`\u8B1B`].string() // U+8B1B <cjk>
	0x76: [`\u8CA2`].string() // U+8CA2 <cjk>
	0x77: [`\u8CFC`].string() // U+8CFC <cjk>
	0x78: [`\u90CA`].string() // U+90CA <cjk>
	0x79: [`\u9175`].string() // U+9175 <cjk>
	0x7A: [`\u9271`].string() // U+9271 <cjk>
	0x7B: [`\u783F`].string() // U+783F <cjk>
	0x7C: [`\u92FC`].string() // U+92FC <cjk>
	0x7D: [`\u95A4`].string() // U+95A4 <cjk>
	0x7E: [`\u964D`].string() // U+964D <cjk>
	0x80: [`\u9805`].string() // U+9805 <cjk>
	0x81: [`\u9999`].string() // U+9999 <cjk>
	0x82: [`\u9AD8`].string() // U+9AD8 <cjk>
	0x83: [`\u9D3B`].string() // U+9D3B <cjk>
	0x84: [`\u525B`].string() // U+525B <cjk>
	0x85: [`\u52AB`].string() // U+52AB <cjk>
	0x86: [`\u53F7`].string() // U+53F7 <cjk>
	0x87: [`\u5408`].string() // U+5408 <cjk>
	0x88: [`\u58D5`].string() // U+58D5 <cjk>
	0x89: [`\u62F7`].string() // U+62F7 <cjk>
	0x8A: [`\u6FE0`].string() // U+6FE0 <cjk>
	0x8B: [`\u8C6A`].string() // U+8C6A <cjk>
	0x8C: [`\u8F5F`].string() // U+8F5F <cjk>
	0x8D: [`\u9EB9`].string() // U+9EB9 <cjk>
	0x8E: [`\u514B`].string() // U+514B <cjk>
	0x8F: [`\u523B`].string() // U+523B <cjk>
	0x90: [`\u544A`].string() // U+544A <cjk>
	0x91: [`\u56FD`].string() // U+56FD <cjk>
	0x92: [`\u7A40`].string() // U+7A40 <cjk>
	0x93: [`\u9177`].string() // U+9177 <cjk>
	0x94: [`\u9D60`].string() // U+9D60 <cjk>
	0x95: [`\u9ED2`].string() // U+9ED2 <cjk>
	0x96: [`\u7344`].string() // U+7344 <cjk>
	0x97: [`\u6F09`].string() // U+6F09 <cjk>
	0x98: [`\u8170`].string() // U+8170 <cjk>
	0x99: [`\u7511`].string() // U+7511 <cjk>
	0x9A: [`\u5FFD`].string() // U+5FFD <cjk>
	0x9B: [`\u60DA`].string() // U+60DA <cjk>
	0x9C: [`\u9AA8`].string() // U+9AA8 <cjk>
	0x9D: [`\u72DB`].string() // U+72DB <cjk>
	0x9E: [`\u8FBC`].string() // U+8FBC <cjk>
	0x9F: [`\u6B64`].string() // U+6B64 <cjk>
	0xA0: [`\u9803`].string() // U+9803 <cjk>
	0xA1: [`\u4ECA`].string() // U+4ECA <cjk>
	0xA2: [`\u56F0`].string() // U+56F0 <cjk>
	0xA3: [`\u5764`].string() // U+5764 <cjk>
	0xA4: [`\u58BE`].string() // U+58BE <cjk>
	0xA5: [`\u5A5A`].string() // U+5A5A <cjk>
	0xA6: [`\u6068`].string() // U+6068 <cjk>
	0xA7: [`\u61C7`].string() // U+61C7 <cjk>
	0xA8: [`\u660F`].string() // U+660F <cjk>
	0xA9: [`\u6606`].string() // U+6606 <cjk>
	0xAA: [`\u6839`].string() // U+6839 <cjk>
	0xAB: [`\u68B1`].string() // U+68B1 <cjk>
	0xAC: [`\u6DF7`].string() // U+6DF7 <cjk>
	0xAD: [`\u75D5`].string() // U+75D5 <cjk>
	0xAE: [`\u7D3A`].string() // U+7D3A <cjk>
	0xAF: [`\u826E`].string() // U+826E <cjk>
	0xB0: [`\u9B42`].string() // U+9B42 <cjk>
	0xB1: [`\u4E9B`].string() // U+4E9B <cjk>
	0xB2: [`\u4F50`].string() // U+4F50 <cjk>
	0xB3: [`\u53C9`].string() // U+53C9 <cjk>
	0xB4: [`\u5506`].string() // U+5506 <cjk>
	0xB5: [`\u5D6F`].string() // U+5D6F <cjk>
	0xB6: [`\u5DE6`].string() // U+5DE6 <cjk>
	0xB7: [`\u5DEE`].string() // U+5DEE <cjk>
	0xB8: [`\u67FB`].string() // U+67FB <cjk>
	0xB9: [`\u6C99`].string() // U+6C99 <cjk>
	0xBA: [`\u7473`].string() // U+7473 <cjk>
	0xBB: [`\u7802`].string() // U+7802 <cjk>
	0xBC: [`\u8A50`].string() // U+8A50 <cjk>
	0xBD: [`\u9396`].string() // U+9396 <cjk>
	0xBE: [`\u88DF`].string() // U+88DF <cjk>
	0xBF: [`\u5750`].string() // U+5750 <cjk>
	0xC0: [`\u5EA7`].string() // U+5EA7 <cjk>
	0xC1: [`\u632B`].string() // U+632B <cjk>
	0xC2: [`\u50B5`].string() // U+50B5 <cjk>
	0xC3: [`\u50AC`].string() // U+50AC <cjk>
	0xC4: [`\u518D`].string() // U+518D <cjk>
	0xC5: [`\u6700`].string() // U+6700 <cjk>
	0xC6: [`\u54C9`].string() // U+54C9 <cjk>
	0xC7: [`\u585E`].string() // U+585E <cjk>
	0xC8: [`\u59BB`].string() // U+59BB <cjk>
	0xC9: [`\u5BB0`].string() // U+5BB0 <cjk>
	0xCA: [`\u5F69`].string() // U+5F69 <cjk>
	0xCB: [`\u624D`].string() // U+624D <cjk>
	0xCC: [`\u63A1`].string() // U+63A1 <cjk>
	0xCD: [`\u683D`].string() // U+683D <cjk>
	0xCE: [`\u6B73`].string() // U+6B73 <cjk>
	0xCF: [`\u6E08`].string() // U+6E08 <cjk>
	0xD0: [`\u707D`].string() // U+707D <cjk>
	0xD1: [`\u91C7`].string() // U+91C7 <cjk>
	0xD2: [`\u7280`].string() // U+7280 <cjk>
	0xD3: [`\u7815`].string() // U+7815 <cjk>
	0xD4: [`\u7826`].string() // U+7826 <cjk>
	0xD5: [`\u796D`].string() // U+796D <cjk>
	0xD6: [`\u658E`].string() // U+658E <cjk>
	0xD7: [`\u7D30`].string() // U+7D30 <cjk>
	0xD8: [`\u83DC`].string() // U+83DC <cjk>
	0xD9: [`\u88C1`].string() // U+88C1 <cjk>
	0xDA: [`\u8F09`].string() // U+8F09 <cjk>
	0xDB: [`\u969B`].string() // U+969B <cjk>
	0xDC: [`\u5264`].string() // U+5264 <cjk>
	0xDD: [`\u5728`].string() // U+5728 <cjk>
	0xDE: [`\u6750`].string() // U+6750 <cjk>
	0xDF: [`\u7F6A`].string() // U+7F6A <cjk>
	0xE0: [`\u8CA1`].string() // U+8CA1 <cjk>
	0xE1: [`\u51B4`].string() // U+51B4 <cjk>
	0xE2: [`\u5742`].string() // U+5742 <cjk>
	0xE3: [`\u962A`].string() // U+962A <cjk>
	0xE4: [`\u583A`].string() // U+583A <cjk>
	0xE5: [`\u698A`].string() // U+698A <cjk>
	0xE6: [`\u80B4`].string() // U+80B4 <cjk>
	0xE7: [`\u54B2`].string() // U+54B2 <cjk>
	0xE8: [`\u5D0E`].string() // U+5D0E <cjk>
	0xE9: [`\u57FC`].string() // U+57FC <cjk>
	0xEA: [`\u7895`].string() // U+7895 <cjk>
	0xEB: [`\u9DFA`].string() // U+9DFA <cjk>
	0xEC: [`\u4F5C`].string() // U+4F5C <cjk>
	0xED: [`\u524A`].string() // U+524A <cjk>
	0xEE: [`\u548B`].string() // U+548B <cjk>
	0xEF: [`\u643E`].string() // U+643E <cjk>
	0xF0: [`\u6628`].string() // U+6628 <cjk>
	0xF1: [`\u6714`].string() // U+6714 <cjk>
	0xF2: [`\u67F5`].string() // U+67F5 <cjk>
	0xF3: [`\u7A84`].string() // U+7A84 <cjk>
	0xF4: [`\u7B56`].string() // U+7B56 <cjk>
	0xF5: [`\u7D22`].string() // U+7D22 <cjk>
	0xF6: [`\u932F`].string() // U+932F <cjk>
	0xF7: [`\u685C`].string() // U+685C <cjk>
	0xF8: [`\u9BAD`].string() // U+9BAD <cjk>
	0xF9: [`\u7B39`].string() // U+7B39 <cjk>
	0xFA: [`\u5319`].string() // U+5319 <cjk>
	0xFB: [`\u518A`].string() // U+518A <cjk>
	0xFC: [`\u5237`].string() // U+5237 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xea = {
	0x40: [`\u9D5D`].string() // U+9D5D <cjk>
	0x41: [`\u9D5E`].string() // U+9D5E <cjk>
	0x42: [`\u9D64`].string() // U+9D64 <cjk>
	0x43: [`\u9D51`].string() // U+9D51 <cjk>
	0x44: [`\u9D50`].string() // U+9D50 <cjk>
	0x45: [`\u9D59`].string() // U+9D59 <cjk>
	0x46: [`\u9D72`].string() // U+9D72 <cjk>
	0x47: [`\u9D89`].string() // U+9D89 <cjk>
	0x48: [`\u9D87`].string() // U+9D87 <cjk>
	0x49: [`\u9DAB`].string() // U+9DAB <cjk>
	0x4A: [`\u9D6F`].string() // U+9D6F <cjk>
	0x4B: [`\u9D7A`].string() // U+9D7A <cjk>
	0x4C: [`\u9D9A`].string() // U+9D9A <cjk>
	0x4D: [`\u9DA4`].string() // U+9DA4 <cjk>
	0x4E: [`\u9DA9`].string() // U+9DA9 <cjk>
	0x4F: [`\u9DB2`].string() // U+9DB2 <cjk>
	0x50: [`\u9DC4`].string() // U+9DC4 <cjk>
	0x51: [`\u9DC1`].string() // U+9DC1 <cjk>
	0x52: [`\u9DBB`].string() // U+9DBB <cjk>
	0x53: [`\u9DB8`].string() // U+9DB8 <cjk>
	0x54: [`\u9DBA`].string() // U+9DBA <cjk>
	0x55: [`\u9DC6`].string() // U+9DC6 <cjk>
	0x56: [`\u9DCF`].string() // U+9DCF <cjk>
	0x57: [`\u9DC2`].string() // U+9DC2 <cjk>
	0x58: [`\u9DD9`].string() // U+9DD9 <cjk>
	0x59: [`\u9DD3`].string() // U+9DD3 <cjk>
	0x5A: [`\u9DF8`].string() // U+9DF8 <cjk>
	0x5B: [`\u9DE6`].string() // U+9DE6 <cjk>
	0x5C: [`\u9DED`].string() // U+9DED <cjk>
	0x5D: [`\u9DEF`].string() // U+9DEF <cjk>
	0x5E: [`\u9DFD`].string() // U+9DFD <cjk>
	0x5F: [`\u9E1A`].string() // U+9E1A <cjk>
	0x60: [`\u9E1B`].string() // U+9E1B <cjk>
	0x61: [`\u9E1E`].string() // U+9E1E <cjk>
	0x62: [`\u9E75`].string() // U+9E75 <cjk>
	0x63: [`\u9E79`].string() // U+9E79 <cjk>
	0x64: [`\u9E7D`].string() // U+9E7D <cjk>
	0x65: [`\u9E81`].string() // U+9E81 <cjk>
	0x66: [`\u9E88`].string() // U+9E88 <cjk>
	0x67: [`\u9E8B`].string() // U+9E8B <cjk>
	0x68: [`\u9E8C`].string() // U+9E8C <cjk>
	0x69: [`\u9E92`].string() // U+9E92 <cjk>
	0x6A: [`\u9E95`].string() // U+9E95 <cjk>
	0x6B: [`\u9E91`].string() // U+9E91 <cjk>
	0x6C: [`\u9E9D`].string() // U+9E9D <cjk>
	0x6D: [`\u9EA5`].string() // U+9EA5 <cjk>
	0x6E: [`\u9EA9`].string() // U+9EA9 <cjk>
	0x6F: [`\u9EB8`].string() // U+9EB8 <cjk>
	0x70: [`\u9EAA`].string() // U+9EAA <cjk>
	0x71: [`\u9EAD`].string() // U+9EAD <cjk>
	0x72: [`\u9761`].string() // U+9761 <cjk>
	0x73: [`\u9ECC`].string() // U+9ECC <cjk>
	0x74: [`\u9ECE`].string() // U+9ECE <cjk>
	0x75: [`\u9ECF`].string() // U+9ECF <cjk>
	0x76: [`\u9ED0`].string() // U+9ED0 <cjk>
	0x77: [`\u9ED4`].string() // U+9ED4 <cjk>
	0x78: [`\u9EDC`].string() // U+9EDC <cjk>
	0x79: [`\u9EDE`].string() // U+9EDE <cjk>
	0x7A: [`\u9EDD`].string() // U+9EDD <cjk>
	0x7B: [`\u9EE0`].string() // U+9EE0 <cjk>
	0x7C: [`\u9EE5`].string() // U+9EE5 <cjk>
	0x7D: [`\u9EE8`].string() // U+9EE8 <cjk>
	0x7E: [`\u9EEF`].string() // U+9EEF <cjk>
	0x80: [`\u9EF4`].string() // U+9EF4 <cjk>
	0x81: [`\u9EF6`].string() // U+9EF6 <cjk>
	0x82: [`\u9EF7`].string() // U+9EF7 <cjk>
	0x83: [`\u9EF9`].string() // U+9EF9 <cjk>
	0x84: [`\u9EFB`].string() // U+9EFB <cjk>
	0x85: [`\u9EFC`].string() // U+9EFC <cjk>
	0x86: [`\u9EFD`].string() // U+9EFD <cjk>
	0x87: [`\u9F07`].string() // U+9F07 <cjk>
	0x88: [`\u9F08`].string() // U+9F08 <cjk>
	0x89: [`\u76B7`].string() // U+76B7 <cjk>
	0x8A: [`\u9F15`].string() // U+9F15 <cjk>
	0x8B: [`\u9F21`].string() // U+9F21 <cjk>
	0x8C: [`\u9F2C`].string() // U+9F2C <cjk>
	0x8D: [`\u9F3E`].string() // U+9F3E <cjk>
	0x8E: [`\u9F4A`].string() // U+9F4A <cjk>
	0x8F: [`\u9F52`].string() // U+9F52 <cjk>
	0x90: [`\u9F54`].string() // U+9F54 <cjk>
	0x91: [`\u9F63`].string() // U+9F63 <cjk>
	0x92: [`\u9F5F`].string() // U+9F5F <cjk>
	0x93: [`\u9F60`].string() // U+9F60 <cjk>
	0x94: [`\u9F61`].string() // U+9F61 <cjk>
	0x95: [`\u9F66`].string() // U+9F66 <cjk>
	0x96: [`\u9F67`].string() // U+9F67 <cjk>
	0x97: [`\u9F6C`].string() // U+9F6C <cjk>
	0x98: [`\u9F6A`].string() // U+9F6A <cjk>
	0x99: [`\u9F77`].string() // U+9F77 <cjk>
	0x9A: [`\u9F72`].string() // U+9F72 <cjk>
	0x9B: [`\u9F76`].string() // U+9F76 <cjk>
	0x9C: [`\u9F95`].string() // U+9F95 <cjk>
	0x9D: [`\u9F9C`].string() // U+9F9C <cjk>
	0x9E: [`\u9FA0`].string() // U+9FA0 <cjk>
	0x9F: [`\u582F`].string() // U+582F <cjk>
	0xA0: [`\u69C7`].string() // U+69C7 <cjk>
	0xA1: [`\u9059`].string() // U+9059 <cjk>
	0xA2: [`\u7464`].string() // U+7464 <cjk>
	0xA3: [`\u51DC`].string() // U+51DC <cjk>
	0xA4: [`\u7199`].string() // U+7199 <cjk>
	0xA5: [`\u5653`].string() // U+5653 <cjk>
	0xA6: [`\u5DE2`].string() // U+5DE2 <cjk>
	0xA7: [`\u5E14`].string() // U+5E14 <cjk>
	0xA8: [`\u5E18`].string() // U+5E18 <cjk>
	0xA9: [`\u5E58`].string() // U+5E58 <cjk>
	0xAA: [`\u5E5E`].string() // U+5E5E <cjk>
	0xAB: [`\u5EBE`].string() // U+5EBE <cjk>
	0xAC: [`\uF928`].string() // U+F928 CJK COMPATIBILITY IDEOGRAPH-F928
	0xAD: [`\u5ECB`].string() // U+5ECB <cjk>
	0xAE: [`\u5EF9`].string() // U+5EF9 <cjk>
	0xAF: [`\u5F00`].string() // U+5F00 <cjk>
	0xB0: [`\u5F02`].string() // U+5F02 <cjk>
	0xB1: [`\u5F07`].string() // U+5F07 <cjk>
	0xB2: [`\u5F1D`].string() // U+5F1D <cjk>
	0xB3: [`\u5F23`].string() // U+5F23 <cjk>
	0xB4: [`\u5F34`].string() // U+5F34 <cjk>
	0xB5: [`\u5F36`].string() // U+5F36 <cjk>
	0xB6: [`\u5F3D`].string() // U+5F3D <cjk>
	0xB7: [`\u5F40`].string() // U+5F40 <cjk>
	0xB8: [`\u5F45`].string() // U+5F45 <cjk>
	0xB9: [`\u5F54`].string() // U+5F54 <cjk>
	0xBA: [`\u5F58`].string() // U+5F58 <cjk>
	0xBB: [`\u5F64`].string() // U+5F64 <cjk>
	0xBC: [`\u5F67`].string() // U+5F67 <cjk>
	0xBD: [`\u5F7D`].string() // U+5F7D <cjk>
	0xBE: [`\u5F89`].string() // U+5F89 <cjk>
	0xBF: [`\u5F9C`].string() // U+5F9C <cjk>
	0xC0: [`\u5FA7`].string() // U+5FA7 <cjk>
	0xC1: [`\u5FAF`].string() // U+5FAF <cjk>
	0xC2: [`\u5FB5`].string() // U+5FB5 <cjk>
	0xC3: [`\u5FB7`].string() // U+5FB7 <cjk>
	0xC4: [`\u5FC9`].string() // U+5FC9 <cjk>
	0xC5: [`\u5FDE`].string() // U+5FDE <cjk>
	0xC6: [`\u5FE1`].string() // U+5FE1 <cjk>
	0xC7: [`\u5FE9`].string() // U+5FE9 <cjk>
	0xC8: [`\u600D`].string() // U+600D <cjk>
	0xC9: [`\u6014`].string() // U+6014 <cjk>
	0xCA: [`\u6018`].string() // U+6018 <cjk>
	0xCB: [`\u6033`].string() // U+6033 <cjk>
	0xCC: [`\u6035`].string() // U+6035 <cjk>
	0xCD: [`\u6047`].string() // U+6047 <cjk>
	0xCE: [`\uFA3D`].string() // U+FA3D CJK COMPATIBILITY IDEOGRAPH-FA3D
	0xCF: [`\u609D`].string() // U+609D <cjk>
	0xD0: [`\u609E`].string() // U+609E <cjk>
	0xD1: [`\u60CB`].string() // U+60CB <cjk>
	0xD2: [`\u60D4`].string() // U+60D4 <cjk>
	0xD3: [`\u60D5`].string() // U+60D5 <cjk>
	0xD4: [`\u60DD`].string() // U+60DD <cjk>
	0xD5: [`\u60F8`].string() // U+60F8 <cjk>
	0xD6: [`\u611C`].string() // U+611C <cjk>
	0xD7: [`\u612B`].string() // U+612B <cjk>
	0xD8: [`\u6130`].string() // U+6130 <cjk>
	0xD9: [`\u6137`].string() // U+6137 <cjk>
	0xDA: [`\uFA3E`].string() // U+FA3E CJK COMPATIBILITY IDEOGRAPH-FA3E
	0xDB: [`\u618D`].string() // U+618D <cjk>
	0xDC: [`\uFA3F`].string() // U+FA3F CJK COMPATIBILITY IDEOGRAPH-FA3F
	0xDD: [`\u61BC`].string() // U+61BC <cjk>
	0xDE: [`\u61B9`].string() // U+61B9 <cjk>
	0xDF: [`\uFA40`].string() // U+FA40 CJK COMPATIBILITY IDEOGRAPH-FA40
	0xE0: [`\u6222`].string() // U+6222 <cjk>
	0xE1: [`\u623E`].string() // U+623E <cjk>
	0xE2: [`\u6243`].string() // U+6243 <cjk>
	0xE3: [`\u6256`].string() // U+6256 <cjk>
	0xE4: [`\u625A`].string() // U+625A <cjk>
	0xE5: [`\u626F`].string() // U+626F <cjk>
	0xE6: [`\u6285`].string() // U+6285 <cjk>
	0xE7: [`\u62C4`].string() // U+62C4 <cjk>
	0xE8: [`\u62D6`].string() // U+62D6 <cjk>
	0xE9: [`\u62FC`].string() // U+62FC <cjk>
	0xEA: [`\u630A`].string() // U+630A <cjk>
	0xEB: [`\u6318`].string() // U+6318 <cjk>
	0xEC: [`\u6339`].string() // U+6339 <cjk>
	0xED: [`\u6343`].string() // U+6343 <cjk>
	0xEE: [`\u6365`].string() // U+6365 <cjk>
	0xEF: [`\u637C`].string() // U+637C <cjk>
	0xF0: [`\u63E5`].string() // U+63E5 <cjk>
	0xF1: [`\u63ED`].string() // U+63ED <cjk>
	0xF2: [`\u63F5`].string() // U+63F5 <cjk>
	0xF3: [`\u6410`].string() // U+6410 <cjk>
	0xF4: [`\u6414`].string() // U+6414 <cjk>
	0xF5: [`\u6422`].string() // U+6422 <cjk>
	0xF6: [`\u6479`].string() // U+6479 <cjk>
	0xF7: [`\u6451`].string() // U+6451 <cjk>
	0xF8: [`\u6460`].string() // U+6460 <cjk>
	0xF9: [`\u646D`].string() // U+646D <cjk>
	0xFA: [`\u64CE`].string() // U+64CE <cjk>
	0xFB: [`\u64BE`].string() // U+64BE <cjk>
	0xFC: [`\u64BF`].string() // U+64BF <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x8a = {
	0x40: [`\u9B41`].string() // U+9B41 <cjk>
	0x41: [`\u6666`].string() // U+6666 <cjk>
	0x42: [`\u68B0`].string() // U+68B0 <cjk>
	0x43: [`\u6D77`].string() // U+6D77 <cjk>
	0x44: [`\u7070`].string() // U+7070 <cjk>
	0x45: [`\u754C`].string() // U+754C <cjk>
	0x46: [`\u7686`].string() // U+7686 <cjk>
	0x47: [`\u7D75`].string() // U+7D75 <cjk>
	0x48: [`\u82A5`].string() // U+82A5 <cjk>
	0x49: [`\u87F9`].string() // U+87F9 <cjk>
	0x4A: [`\u958B`].string() // U+958B <cjk>
	0x4B: [`\u968E`].string() // U+968E <cjk>
	0x4C: [`\u8C9D`].string() // U+8C9D <cjk>
	0x4D: [`\u51F1`].string() // U+51F1 <cjk>
	0x4E: [`\u52BE`].string() // U+52BE <cjk>
	0x4F: [`\u5916`].string() // U+5916 <cjk>
	0x50: [`\u54B3`].string() // U+54B3 <cjk>
	0x51: [`\u5BB3`].string() // U+5BB3 <cjk>
	0x52: [`\u5D16`].string() // U+5D16 <cjk>
	0x53: [`\u6168`].string() // U+6168 <cjk>
	0x54: [`\u6982`].string() // U+6982 <cjk>
	0x55: [`\u6DAF`].string() // U+6DAF <cjk>
	0x56: [`\u788D`].string() // U+788D <cjk>
	0x57: [`\u84CB`].string() // U+84CB <cjk>
	0x58: [`\u8857`].string() // U+8857 <cjk>
	0x59: [`\u8A72`].string() // U+8A72 <cjk>
	0x5A: [`\u93A7`].string() // U+93A7 <cjk>
	0x5B: [`\u9AB8`].string() // U+9AB8 <cjk>
	0x5C: [`\u6D6C`].string() // U+6D6C <cjk>
	0x5D: [`\u99A8`].string() // U+99A8 <cjk>
	0x5E: [`\u86D9`].string() // U+86D9 <cjk>
	0x5F: [`\u57A3`].string() // U+57A3 <cjk>
	0x60: [`\u67FF`].string() // U+67FF <cjk>
	0x61: [`\u86CE`].string() // U+86CE <cjk>
	0x62: [`\u920E`].string() // U+920E <cjk>
	0x63: [`\u5283`].string() // U+5283 <cjk>
	0x64: [`\u5687`].string() // U+5687 <cjk>
	0x65: [`\u5404`].string() // U+5404 <cjk>
	0x66: [`\u5ED3`].string() // U+5ED3 <cjk>
	0x67: [`\u62E1`].string() // U+62E1 <cjk>
	0x68: [`\u64B9`].string() // U+64B9 <cjk>
	0x69: [`\u683C`].string() // U+683C <cjk>
	0x6A: [`\u6838`].string() // U+6838 <cjk>
	0x6B: [`\u6BBB`].string() // U+6BBB <cjk>
	0x6C: [`\u7372`].string() // U+7372 <cjk>
	0x6D: [`\u78BA`].string() // U+78BA <cjk>
	0x6E: [`\u7A6B`].string() // U+7A6B <cjk>
	0x6F: [`\u899A`].string() // U+899A <cjk>
	0x70: [`\u89D2`].string() // U+89D2 <cjk>
	0x71: [`\u8D6B`].string() // U+8D6B <cjk>
	0x72: [`\u8F03`].string() // U+8F03 <cjk>
	0x73: [`\u90ED`].string() // U+90ED <cjk>
	0x74: [`\u95A3`].string() // U+95A3 <cjk>
	0x75: [`\u9694`].string() // U+9694 <cjk>
	0x76: [`\u9769`].string() // U+9769 <cjk>
	0x77: [`\u5B66`].string() // U+5B66 <cjk>
	0x78: [`\u5CB3`].string() // U+5CB3 <cjk>
	0x79: [`\u697D`].string() // U+697D <cjk>
	0x7A: [`\u984D`].string() // U+984D <cjk>
	0x7B: [`\u984E`].string() // U+984E <cjk>
	0x7C: [`\u639B`].string() // U+639B <cjk>
	0x7D: [`\u7B20`].string() // U+7B20 <cjk>
	0x7E: [`\u6A2B`].string() // U+6A2B <cjk>
	0x80: [`\u6A7F`].string() // U+6A7F <cjk>
	0x81: [`\u68B6`].string() // U+68B6 <cjk>
	0x82: [`\u9C0D`].string() // U+9C0D <cjk>
	0x83: [`\u6F5F`].string() // U+6F5F <cjk>
	0x84: [`\u5272`].string() // U+5272 <cjk>
	0x85: [`\u559D`].string() // U+559D <cjk>
	0x86: [`\u6070`].string() // U+6070 <cjk>
	0x87: [`\u62EC`].string() // U+62EC <cjk>
	0x88: [`\u6D3B`].string() // U+6D3B <cjk>
	0x89: [`\u6E07`].string() // U+6E07 <cjk>
	0x8A: [`\u6ED1`].string() // U+6ED1 <cjk>
	0x8B: [`\u845B`].string() // U+845B <cjk>
	0x8C: [`\u8910`].string() // U+8910 <cjk>
	0x8D: [`\u8F44`].string() // U+8F44 <cjk>
	0x8E: [`\u4E14`].string() // U+4E14 <cjk>
	0x8F: [`\u9C39`].string() // U+9C39 <cjk>
	0x90: [`\u53F6`].string() // U+53F6 <cjk>
	0x91: [`\u691B`].string() // U+691B <cjk>
	0x92: [`\u6A3A`].string() // U+6A3A <cjk>
	0x93: [`\u9784`].string() // U+9784 <cjk>
	0x94: [`\u682A`].string() // U+682A <cjk>
	0x95: [`\u515C`].string() // U+515C <cjk>
	0x96: [`\u7AC3`].string() // U+7AC3 <cjk>
	0x97: [`\u84B2`].string() // U+84B2 <cjk>
	0x98: [`\u91DC`].string() // U+91DC <cjk>
	0x99: [`\u938C`].string() // U+938C <cjk>
	0x9A: [`\u565B`].string() // U+565B <cjk>
	0x9B: [`\u9D28`].string() // U+9D28 <cjk>
	0x9C: [`\u6822`].string() // U+6822 <cjk>
	0x9D: [`\u8305`].string() // U+8305 <cjk>
	0x9E: [`\u8431`].string() // U+8431 <cjk>
	0x9F: [`\u7CA5`].string() // U+7CA5 <cjk>
	0xA0: [`\u5208`].string() // U+5208 <cjk>
	0xA1: [`\u82C5`].string() // U+82C5 <cjk>
	0xA2: [`\u74E6`].string() // U+74E6 <cjk>
	0xA3: [`\u4E7E`].string() // U+4E7E <cjk>
	0xA4: [`\u4F83`].string() // U+4F83 <cjk>
	0xA5: [`\u51A0`].string() // U+51A0 <cjk>
	0xA6: [`\u5BD2`].string() // U+5BD2 <cjk>
	0xA7: [`\u520A`].string() // U+520A <cjk>
	0xA8: [`\u52D8`].string() // U+52D8 <cjk>
	0xA9: [`\u52E7`].string() // U+52E7 <cjk>
	0xAA: [`\u5DFB`].string() // U+5DFB <cjk>
	0xAB: [`\u559A`].string() // U+559A <cjk>
	0xAC: [`\u582A`].string() // U+582A <cjk>
	0xAD: [`\u59E6`].string() // U+59E6 <cjk>
	0xAE: [`\u5B8C`].string() // U+5B8C <cjk>
	0xAF: [`\u5B98`].string() // U+5B98 <cjk>
	0xB0: [`\u5BDB`].string() // U+5BDB <cjk>
	0xB1: [`\u5E72`].string() // U+5E72 <cjk>
	0xB2: [`\u5E79`].string() // U+5E79 <cjk>
	0xB3: [`\u60A3`].string() // U+60A3 <cjk>
	0xB4: [`\u611F`].string() // U+611F <cjk>
	0xB5: [`\u6163`].string() // U+6163 <cjk>
	0xB6: [`\u61BE`].string() // U+61BE <cjk>
	0xB7: [`\u63DB`].string() // U+63DB <cjk>
	0xB8: [`\u6562`].string() // U+6562 <cjk>
	0xB9: [`\u67D1`].string() // U+67D1 <cjk>
	0xBA: [`\u6853`].string() // U+6853 <cjk>
	0xBB: [`\u68FA`].string() // U+68FA <cjk>
	0xBC: [`\u6B3E`].string() // U+6B3E <cjk>
	0xBD: [`\u6B53`].string() // U+6B53 <cjk>
	0xBE: [`\u6C57`].string() // U+6C57 <cjk>
	0xBF: [`\u6F22`].string() // U+6F22 <cjk>
	0xC0: [`\u6F97`].string() // U+6F97 <cjk>
	0xC1: [`\u6F45`].string() // U+6F45 <cjk>
	0xC2: [`\u74B0`].string() // U+74B0 <cjk>
	0xC3: [`\u7518`].string() // U+7518 <cjk>
	0xC4: [`\u76E3`].string() // U+76E3 <cjk>
	0xC5: [`\u770B`].string() // U+770B <cjk>
	0xC6: [`\u7AFF`].string() // U+7AFF <cjk>
	0xC7: [`\u7BA1`].string() // U+7BA1 <cjk>
	0xC8: [`\u7C21`].string() // U+7C21 <cjk>
	0xC9: [`\u7DE9`].string() // U+7DE9 <cjk>
	0xCA: [`\u7F36`].string() // U+7F36 <cjk>
	0xCB: [`\u7FF0`].string() // U+7FF0 <cjk>
	0xCC: [`\u809D`].string() // U+809D <cjk>
	0xCD: [`\u8266`].string() // U+8266 <cjk>
	0xCE: [`\u839E`].string() // U+839E <cjk>
	0xCF: [`\u89B3`].string() // U+89B3 <cjk>
	0xD0: [`\u8ACC`].string() // U+8ACC <cjk>
	0xD1: [`\u8CAB`].string() // U+8CAB <cjk>
	0xD2: [`\u9084`].string() // U+9084 <cjk>
	0xD3: [`\u9451`].string() // U+9451 <cjk>
	0xD4: [`\u9593`].string() // U+9593 <cjk>
	0xD5: [`\u9591`].string() // U+9591 <cjk>
	0xD6: [`\u95A2`].string() // U+95A2 <cjk>
	0xD7: [`\u9665`].string() // U+9665 <cjk>
	0xD8: [`\u97D3`].string() // U+97D3 <cjk>
	0xD9: [`\u9928`].string() // U+9928 <cjk>
	0xDA: [`\u8218`].string() // U+8218 <cjk>
	0xDB: [`\u4E38`].string() // U+4E38 <cjk>
	0xDC: [`\u542B`].string() // U+542B <cjk>
	0xDD: [`\u5CB8`].string() // U+5CB8 <cjk>
	0xDE: [`\u5DCC`].string() // U+5DCC <cjk>
	0xDF: [`\u73A9`].string() // U+73A9 <cjk>
	0xE0: [`\u764C`].string() // U+764C <cjk>
	0xE1: [`\u773C`].string() // U+773C <cjk>
	0xE2: [`\u5CA9`].string() // U+5CA9 <cjk>
	0xE3: [`\u7FEB`].string() // U+7FEB <cjk>
	0xE4: [`\u8D0B`].string() // U+8D0B <cjk>
	0xE5: [`\u96C1`].string() // U+96C1 <cjk>
	0xE6: [`\u9811`].string() // U+9811 <cjk>
	0xE7: [`\u9854`].string() // U+9854 <cjk>
	0xE8: [`\u9858`].string() // U+9858 <cjk>
	0xE9: [`\u4F01`].string() // U+4F01 <cjk>
	0xEA: [`\u4F0E`].string() // U+4F0E <cjk>
	0xEB: [`\u5371`].string() // U+5371 <cjk>
	0xEC: [`\u559C`].string() // U+559C <cjk>
	0xED: [`\u5668`].string() // U+5668 <cjk>
	0xEE: [`\u57FA`].string() // U+57FA <cjk>
	0xEF: [`\u5947`].string() // U+5947 <cjk>
	0xF0: [`\u5B09`].string() // U+5B09 <cjk>
	0xF1: [`\u5BC4`].string() // U+5BC4 <cjk>
	0xF2: [`\u5C90`].string() // U+5C90 <cjk>
	0xF3: [`\u5E0C`].string() // U+5E0C <cjk>
	0xF4: [`\u5E7E`].string() // U+5E7E <cjk>
	0xF5: [`\u5FCC`].string() // U+5FCC <cjk>
	0xF6: [`\u63EE`].string() // U+63EE <cjk>
	0xF7: [`\u673A`].string() // U+673A <cjk>
	0xF8: [`\u65D7`].string() // U+65D7 <cjk>
	0xF9: [`\u65E2`].string() // U+65E2 <cjk>
	0xFA: [`\u671F`].string() // U+671F <cjk>
	0xFB: [`\u68CB`].string() // U+68CB <cjk>
	0xFC: [`\u68C4`].string() // U+68C4 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x9b = {
	0x40: [`\u5978`].string() // U+5978 <cjk>
	0x41: [`\u5981`].string() // U+5981 <cjk>
	0x42: [`\u599D`].string() // U+599D <cjk>
	0x43: [`\u4F5E`].string() // U+4F5E <cjk>
	0x44: [`\u4FAB`].string() // U+4FAB <cjk>
	0x45: [`\u59A3`].string() // U+59A3 <cjk>
	0x46: [`\u59B2`].string() // U+59B2 <cjk>
	0x47: [`\u59C6`].string() // U+59C6 <cjk>
	0x48: [`\u59E8`].string() // U+59E8 <cjk>
	0x49: [`\u59DC`].string() // U+59DC <cjk>
	0x4A: [`\u598D`].string() // U+598D <cjk>
	0x4B: [`\u59D9`].string() // U+59D9 <cjk>
	0x4C: [`\u59DA`].string() // U+59DA <cjk>
	0x4D: [`\u5A25`].string() // U+5A25 <cjk>
	0x4E: [`\u5A1F`].string() // U+5A1F <cjk>
	0x4F: [`\u5A11`].string() // U+5A11 <cjk>
	0x50: [`\u5A1C`].string() // U+5A1C <cjk>
	0x51: [`\u5A09`].string() // U+5A09 <cjk>
	0x52: [`\u5A1A`].string() // U+5A1A <cjk>
	0x53: [`\u5A40`].string() // U+5A40 <cjk>
	0x54: [`\u5A6C`].string() // U+5A6C <cjk>
	0x55: [`\u5A49`].string() // U+5A49 <cjk>
	0x56: [`\u5A35`].string() // U+5A35 <cjk>
	0x57: [`\u5A36`].string() // U+5A36 <cjk>
	0x58: [`\u5A62`].string() // U+5A62 <cjk>
	0x59: [`\u5A6A`].string() // U+5A6A <cjk>
	0x5A: [`\u5A9A`].string() // U+5A9A <cjk>
	0x5B: [`\u5ABC`].string() // U+5ABC <cjk>
	0x5C: [`\u5ABE`].string() // U+5ABE <cjk>
	0x5D: [`\u5ACB`].string() // U+5ACB <cjk>
	0x5E: [`\u5AC2`].string() // U+5AC2 <cjk>
	0x5F: [`\u5ABD`].string() // U+5ABD <cjk>
	0x60: [`\u5AE3`].string() // U+5AE3 <cjk>
	0x61: [`\u5AD7`].string() // U+5AD7 <cjk>
	0x62: [`\u5AE6`].string() // U+5AE6 <cjk>
	0x63: [`\u5AE9`].string() // U+5AE9 <cjk>
	0x64: [`\u5AD6`].string() // U+5AD6 <cjk>
	0x65: [`\u5AFA`].string() // U+5AFA <cjk>
	0x66: [`\u5AFB`].string() // U+5AFB <cjk>
	0x67: [`\u5B0C`].string() // U+5B0C <cjk>
	0x68: [`\u5B0B`].string() // U+5B0B <cjk>
	0x69: [`\u5B16`].string() // U+5B16 <cjk>
	0x6A: [`\u5B32`].string() // U+5B32 <cjk>
	0x6B: [`\u5AD0`].string() // U+5AD0 <cjk>
	0x6C: [`\u5B2A`].string() // U+5B2A <cjk>
	0x6D: [`\u5B36`].string() // U+5B36 <cjk>
	0x6E: [`\u5B3E`].string() // U+5B3E <cjk>
	0x6F: [`\u5B43`].string() // U+5B43 <cjk>
	0x70: [`\u5B45`].string() // U+5B45 <cjk>
	0x71: [`\u5B40`].string() // U+5B40 <cjk>
	0x72: [`\u5B51`].string() // U+5B51 <cjk>
	0x73: [`\u5B55`].string() // U+5B55 <cjk>
	0x74: [`\u5B5A`].string() // U+5B5A <cjk>
	0x75: [`\u5B5B`].string() // U+5B5B <cjk>
	0x76: [`\u5B65`].string() // U+5B65 <cjk>
	0x77: [`\u5B69`].string() // U+5B69 <cjk>
	0x78: [`\u5B70`].string() // U+5B70 <cjk>
	0x79: [`\u5B73`].string() // U+5B73 <cjk>
	0x7A: [`\u5B75`].string() // U+5B75 <cjk>
	0x7B: [`\u5B78`].string() // U+5B78 <cjk>
	0x7C: [`\u6588`].string() // U+6588 <cjk>
	0x7D: [`\u5B7A`].string() // U+5B7A <cjk>
	0x7E: [`\u5B80`].string() // U+5B80 <cjk>
	0x80: [`\u5B83`].string() // U+5B83 <cjk>
	0x81: [`\u5BA6`].string() // U+5BA6 <cjk>
	0x82: [`\u5BB8`].string() // U+5BB8 <cjk>
	0x83: [`\u5BC3`].string() // U+5BC3 <cjk>
	0x84: [`\u5BC7`].string() // U+5BC7 <cjk>
	0x85: [`\u5BC9`].string() // U+5BC9 <cjk>
	0x86: [`\u5BD4`].string() // U+5BD4 <cjk>
	0x87: [`\u5BD0`].string() // U+5BD0 <cjk>
	0x88: [`\u5BE4`].string() // U+5BE4 <cjk>
	0x89: [`\u5BE6`].string() // U+5BE6 <cjk>
	0x8A: [`\u5BE2`].string() // U+5BE2 <cjk>
	0x8B: [`\u5BDE`].string() // U+5BDE <cjk>
	0x8C: [`\u5BE5`].string() // U+5BE5 <cjk>
	0x8D: [`\u5BEB`].string() // U+5BEB <cjk>
	0x8E: [`\u5BF0`].string() // U+5BF0 <cjk>
	0x8F: [`\u5BF6`].string() // U+5BF6 <cjk>
	0x90: [`\u5BF3`].string() // U+5BF3 <cjk>
	0x91: [`\u5C05`].string() // U+5C05 <cjk>
	0x92: [`\u5C07`].string() // U+5C07 <cjk>
	0x93: [`\u5C08`].string() // U+5C08 <cjk>
	0x94: [`\u5C0D`].string() // U+5C0D <cjk>
	0x95: [`\u5C13`].string() // U+5C13 <cjk>
	0x96: [`\u5C20`].string() // U+5C20 <cjk>
	0x97: [`\u5C22`].string() // U+5C22 <cjk>
	0x98: [`\u5C28`].string() // U+5C28 <cjk>
	0x99: [`\u5C38`].string() // U+5C38 <cjk>
	0x9A: [`\u5C39`].string() // U+5C39 <cjk>
	0x9B: [`\u5C41`].string() // U+5C41 <cjk>
	0x9C: [`\u5C46`].string() // U+5C46 <cjk>
	0x9D: [`\u5C4E`].string() // U+5C4E <cjk>
	0x9E: [`\u5C53`].string() // U+5C53 <cjk>
	0x9F: [`\u5C50`].string() // U+5C50 <cjk>
	0xA0: [`\u5C4F`].string() // U+5C4F <cjk>
	0xA1: [`\u5B71`].string() // U+5B71 <cjk>
	0xA2: [`\u5C6C`].string() // U+5C6C <cjk>
	0xA3: [`\u5C6E`].string() // U+5C6E <cjk>
	0xA4: [`\u4E62`].string() // U+4E62 <cjk>
	0xA5: [`\u5C76`].string() // U+5C76 <cjk>
	0xA6: [`\u5C79`].string() // U+5C79 <cjk>
	0xA7: [`\u5C8C`].string() // U+5C8C <cjk>
	0xA8: [`\u5C91`].string() // U+5C91 <cjk>
	0xA9: [`\u5C94`].string() // U+5C94 <cjk>
	0xAA: [`\u599B`].string() // U+599B <cjk>
	0xAB: [`\u5CAB`].string() // U+5CAB <cjk>
	0xAC: [`\u5CBB`].string() // U+5CBB <cjk>
	0xAD: [`\u5CB6`].string() // U+5CB6 <cjk>
	0xAE: [`\u5CBC`].string() // U+5CBC <cjk>
	0xAF: [`\u5CB7`].string() // U+5CB7 <cjk>
	0xB0: [`\u5CC5`].string() // U+5CC5 <cjk>
	0xB1: [`\u5CBE`].string() // U+5CBE <cjk>
	0xB2: [`\u5CC7`].string() // U+5CC7 <cjk>
	0xB3: [`\u5CD9`].string() // U+5CD9 <cjk>
	0xB4: [`\u5CE9`].string() // U+5CE9 <cjk>
	0xB5: [`\u5CFD`].string() // U+5CFD <cjk>
	0xB6: [`\u5CFA`].string() // U+5CFA <cjk>
	0xB7: [`\u5CED`].string() // U+5CED <cjk>
	0xB8: [`\u5D8C`].string() // U+5D8C <cjk>
	0xB9: [`\u5CEA`].string() // U+5CEA <cjk>
	0xBA: [`\u5D0B`].string() // U+5D0B <cjk>
	0xBB: [`\u5D15`].string() // U+5D15 <cjk>
	0xBC: [`\u5D17`].string() // U+5D17 <cjk>
	0xBD: [`\u5D5C`].string() // U+5D5C <cjk>
	0xBE: [`\u5D1F`].string() // U+5D1F <cjk>
	0xBF: [`\u5D1B`].string() // U+5D1B <cjk>
	0xC0: [`\u5D11`].string() // U+5D11 <cjk>
	0xC1: [`\u5D14`].string() // U+5D14 <cjk>
	0xC2: [`\u5D22`].string() // U+5D22 <cjk>
	0xC3: [`\u5D1A`].string() // U+5D1A <cjk>
	0xC4: [`\u5D19`].string() // U+5D19 <cjk>
	0xC5: [`\u5D18`].string() // U+5D18 <cjk>
	0xC6: [`\u5D4C`].string() // U+5D4C <cjk>
	0xC7: [`\u5D52`].string() // U+5D52 <cjk>
	0xC8: [`\u5D4E`].string() // U+5D4E <cjk>
	0xC9: [`\u5D4B`].string() // U+5D4B <cjk>
	0xCA: [`\u5D6C`].string() // U+5D6C <cjk>
	0xCB: [`\u5D73`].string() // U+5D73 <cjk>
	0xCC: [`\u5D76`].string() // U+5D76 <cjk>
	0xCD: [`\u5D87`].string() // U+5D87 <cjk>
	0xCE: [`\u5D84`].string() // U+5D84 <cjk>
	0xCF: [`\u5D82`].string() // U+5D82 <cjk>
	0xD0: [`\u5DA2`].string() // U+5DA2 <cjk>
	0xD1: [`\u5D9D`].string() // U+5D9D <cjk>
	0xD2: [`\u5DAC`].string() // U+5DAC <cjk>
	0xD3: [`\u5DAE`].string() // U+5DAE <cjk>
	0xD4: [`\u5DBD`].string() // U+5DBD <cjk>
	0xD5: [`\u5D90`].string() // U+5D90 <cjk>
	0xD6: [`\u5DB7`].string() // U+5DB7 <cjk>
	0xD7: [`\u5DBC`].string() // U+5DBC <cjk>
	0xD8: [`\u5DC9`].string() // U+5DC9 <cjk>
	0xD9: [`\u5DCD`].string() // U+5DCD <cjk>
	0xDA: [`\u5DD3`].string() // U+5DD3 <cjk>
	0xDB: [`\u5DD2`].string() // U+5DD2 <cjk>
	0xDC: [`\u5DD6`].string() // U+5DD6 <cjk>
	0xDD: [`\u5DDB`].string() // U+5DDB <cjk>
	0xDE: [`\u5DEB`].string() // U+5DEB <cjk>
	0xDF: [`\u5DF2`].string() // U+5DF2 <cjk>
	0xE0: [`\u5DF5`].string() // U+5DF5 <cjk>
	0xE1: [`\u5E0B`].string() // U+5E0B <cjk>
	0xE2: [`\u5E1A`].string() // U+5E1A <cjk>
	0xE3: [`\u5E19`].string() // U+5E19 <cjk>
	0xE4: [`\u5E11`].string() // U+5E11 <cjk>
	0xE5: [`\u5E1B`].string() // U+5E1B <cjk>
	0xE6: [`\u5E36`].string() // U+5E36 <cjk>
	0xE7: [`\u5E37`].string() // U+5E37 <cjk>
	0xE8: [`\u5E44`].string() // U+5E44 <cjk>
	0xE9: [`\u5E43`].string() // U+5E43 <cjk>
	0xEA: [`\u5E40`].string() // U+5E40 <cjk>
	0xEB: [`\u5E4E`].string() // U+5E4E <cjk>
	0xEC: [`\u5E57`].string() // U+5E57 <cjk>
	0xED: [`\u5E54`].string() // U+5E54 <cjk>
	0xEE: [`\u5E5F`].string() // U+5E5F <cjk>
	0xEF: [`\u5E62`].string() // U+5E62 <cjk>
	0xF0: [`\u5E64`].string() // U+5E64 <cjk>
	0xF1: [`\u5E47`].string() // U+5E47 <cjk>
	0xF2: [`\u5E75`].string() // U+5E75 <cjk>
	0xF3: [`\u5E76`].string() // U+5E76 <cjk>
	0xF4: [`\u5E7A`].string() // U+5E7A <cjk>
	0xF5: [`\u9EBC`].string() // U+9EBC <cjk>
	0xF6: [`\u5E7F`].string() // U+5E7F <cjk>
	0xF7: [`\u5EA0`].string() // U+5EA0 <cjk>
	0xF8: [`\u5EC1`].string() // U+5EC1 <cjk>
	0xF9: [`\u5EC2`].string() // U+5EC2 <cjk>
	0xFA: [`\u5EC8`].string() // U+5EC8 <cjk>
	0xFB: [`\u5ED0`].string() // U+5ED0 <cjk>
	0xFC: [`\u5ECF`].string() // U+5ECF <cjk>
}

module mojibake

const jis_x_0213_to_utf8_data = {
	0x5C: '¥' // U+00A5 YEN SIGN
	0x7E: '‾' // U+203E OVERLINE
	0xA1: '｡' // U+FF61 HALFWIDTH IDEOGRAPHIC FULL STOP
	0xA2: '｢' // U+FF62 HALFWIDTH LEFT CORNER BRACKET
	0xA3: '｣' // U+FF63 HALFWIDTH RIGHT CORNER BRACKET
	0xA4: '､' // U+FF64 HALFWIDTH IDEOGRAPHIC COMMA
	0xA5: '･' // U+FF65 HALFWIDTH KATAKANA MIDDLE DOT
	0xA6: 'ｦ' // U+FF66 HALFWIDTH KATAKANA LETTER WO
	0xA7: 'ｧ' // U+FF67 HALFWIDTH KATAKANA LETTER SMALL A
	0xA8: 'ｨ' // U+FF68 HALFWIDTH KATAKANA LETTER SMALL I
	0xA9: 'ｩ' // U+FF69 HALFWIDTH KATAKANA LETTER SMALL U
	0xAA: 'ｪ' // U+FF6A HALFWIDTH KATAKANA LETTER SMALL E
	0xAB: 'ｫ' // U+FF6B HALFWIDTH KATAKANA LETTER SMALL O
	0xAC: 'ｬ' // U+FF6C HALFWIDTH KATAKANA LETTER SMALL YA
	0xAD: 'ｭ' // U+FF6D HALFWIDTH KATAKANA LETTER SMALL YU
	0xAE: 'ｮ' // U+FF6E HALFWIDTH KATAKANA LETTER SMALL YO
	0xAF: 'ｯ' // U+FF6F HALFWIDTH KATAKANA LETTER SMALL TU
	0xB0: 'ｰ' // U+FF70 HALFWIDTH KATAKANA-HIRAGANA PROLONGED SOUND MARK
	0xB1: 'ｱ' // U+FF71 HALFWIDTH KATAKANA LETTER A
	0xB2: 'ｲ' // U+FF72 HALFWIDTH KATAKANA LETTER I
	0xB3: 'ｳ' // U+FF73 HALFWIDTH KATAKANA LETTER U
	0xB4: 'ｴ' // U+FF74 HALFWIDTH KATAKANA LETTER E
	0xB5: 'ｵ' // U+FF75 HALFWIDTH KATAKANA LETTER O
	0xB6: 'ｶ' // U+FF76 HALFWIDTH KATAKANA LETTER KA
	0xB7: 'ｷ' // U+FF77 HALFWIDTH KATAKANA LETTER KI
	0xB8: 'ｸ' // U+FF78 HALFWIDTH KATAKANA LETTER KU
	0xB9: 'ｹ' // U+FF79 HALFWIDTH KATAKANA LETTER KE
	0xBA: 'ｺ' // U+FF7A HALFWIDTH KATAKANA LETTER KO
	0xBB: 'ｻ' // U+FF7B HALFWIDTH KATAKANA LETTER SA
	0xBC: 'ｼ' // U+FF7C HALFWIDTH KATAKANA LETTER SI
	0xBD: 'ｽ' // U+FF7D HALFWIDTH KATAKANA LETTER SU
	0xBE: 'ｾ' // U+FF7E HALFWIDTH KATAKANA LETTER SE
	0xBF: 'ｿ' // U+FF7F HALFWIDTH KATAKANA LETTER SO
	0xC0: 'ﾀ' // U+FF80 HALFWIDTH KATAKANA LETTER TA
	0xC1: 'ﾁ' // U+FF81 HALFWIDTH KATAKANA LETTER TI
	0xC2: 'ﾂ' // U+FF82 HALFWIDTH KATAKANA LETTER TU
	0xC3: 'ﾃ' // U+FF83 HALFWIDTH KATAKANA LETTER TE
	0xC4: 'ﾄ' // U+FF84 HALFWIDTH KATAKANA LETTER TO
	0xC5: 'ﾅ' // U+FF85 HALFWIDTH KATAKANA LETTER NA
	0xC6: 'ﾆ' // U+FF86 HALFWIDTH KATAKANA LETTER NI
	0xC7: 'ﾇ' // U+FF87 HALFWIDTH KATAKANA LETTER NU
	0xC8: 'ﾈ' // U+FF88 HALFWIDTH KATAKANA LETTER NE
	0xC9: 'ﾉ' // U+FF89 HALFWIDTH KATAKANA LETTER NO
	0xCA: 'ﾊ' // U+FF8A HALFWIDTH KATAKANA LETTER HA
	0xCB: 'ﾋ' // U+FF8B HALFWIDTH KATAKANA LETTER HI
	0xCC: 'ﾌ' // U+FF8C HALFWIDTH KATAKANA LETTER HU
	0xCD: 'ﾍ' // U+FF8D HALFWIDTH KATAKANA LETTER HE
	0xCE: 'ﾎ' // U+FF8E HALFWIDTH KATAKANA LETTER HO
	0xCF: 'ﾏ' // U+FF8F HALFWIDTH KATAKANA LETTER MA
	0xD0: 'ﾐ' // U+FF90 HALFWIDTH KATAKANA LETTER MI
	0xD1: 'ﾑ' // U+FF91 HALFWIDTH KATAKANA LETTER MU
	0xD2: 'ﾒ' // U+FF92 HALFWIDTH KATAKANA LETTER ME
	0xD3: 'ﾓ' // U+FF93 HALFWIDTH KATAKANA LETTER MO
	0xD4: 'ﾔ' // U+FF94 HALFWIDTH KATAKANA LETTER YA
	0xD5: 'ﾕ' // U+FF95 HALFWIDTH KATAKANA LETTER YU
	0xD6: 'ﾖ' // U+FF96 HALFWIDTH KATAKANA LETTER YO
	0xD7: 'ﾗ' // U+FF97 HALFWIDTH KATAKANA LETTER RA
	0xD8: 'ﾘ' // U+FF98 HALFWIDTH KATAKANA LETTER RI
	0xD9: 'ﾙ' // U+FF99 HALFWIDTH KATAKANA LETTER RU
	0xDA: 'ﾚ' // U+FF9A HALFWIDTH KATAKANA LETTER RE
	0xDB: 'ﾛ' // U+FF9B HALFWIDTH KATAKANA LETTER RO
	0xDC: 'ﾜ' // U+FF9C HALFWIDTH KATAKANA LETTER WA
	0xDD: 'ﾝ' // U+FF9D HALFWIDTH KATAKANA LETTER N
	0xDE: 'ﾞ' // U+FF9E HALFWIDTH KATAKANA VOICED SOUND MARK
	0xDF: 'ﾟ' // U+FF9F HALFWIDTH KATAKANA SEMI-VOICED SOUND MARK
	0x8140: '　' // U+3000 IDEOGRAPHIC SPACE
	0x8141: '、' // U+3001 IDEOGRAPHIC COMMA
	0x8142: '。' // U+3002 IDEOGRAPHIC FULL STOP
	0x8143: '，' // U+FF0C FULLWIDTH COMMA
	0x8144: '．' // U+FF0E FULLWIDTH FULL STOP
	0x8145: '・' // U+30FB KATAKANA MIDDLE DOT
	0x8146: '：' // U+FF1A FULLWIDTH COLON
	0x8147: '；' // U+FF1B FULLWIDTH SEMICOLON
	0x8148: '？' // U+FF1F FULLWIDTH QUESTION MARK
	0x8149: '！' // U+FF01 FULLWIDTH EXCLAMATION MARK
	0x814A: '゛' // U+309B KATAKANA-HIRAGANA VOICED SOUND MARK
	0x814B: '゜' // U+309C KATAKANA-HIRAGANA SEMI-VOICED SOUND MARK
	0x814C: '´' // U+00B4 ACUTE ACCENT
	0x814D: '｀' // U+FF40 FULLWIDTH GRAVE ACCENT
	0x814E: '¨' // U+00A8 DIAERESIS
	0x814F: '＾' // U+FF3E FULLWIDTH CIRCUMFLEX ACCENT
	0x8150: '￣' // U+FFE3 FULLWIDTH MACRON
	0x8151: '＿' // U+FF3F FULLWIDTH LOW LINE
	0x8152: 'ヽ' // U+30FD KATAKANA ITERATION MARK
	0x8153: 'ヾ' // U+30FE KATAKANA VOICED ITERATION MARK
	0x8154: 'ゝ' // U+309D HIRAGANA ITERATION MARK
	0x8155: 'ゞ' // U+309E HIRAGANA VOICED ITERATION MARK
	0x8156: '〃' // U+3003 DITTO MARK
	0x8157: '仝' // U+4EDD <cjk>
	0x8158: '々' // U+3005 IDEOGRAPHIC ITERATION MARK
	0x8159: '〆' // U+3006 IDEOGRAPHIC CLOSING MARK
	0x815A: '〇' // U+3007 IDEOGRAPHIC NUMBER ZERO
	0x815B: 'ー' // U+30FC KATAKANA-HIRAGANA PROLONGED SOUND MARK
	0x815C: '—' // U+2014 EM DASH
	0x815D: '‐' // U+2010 HYPHEN
	0x815E: '／' // U+FF0F FULLWIDTH SOLIDUS
	0x815F: '\\' // U+005C REVERSE SOLIDUS
	0x8160: '〜' // U+301C WAVE DASH
	0x8161: '‖' // U+2016 DOUBLE VERTICAL LINE
	0x8162: '｜' // U+FF5C FULLWIDTH VERTICAL LINE
	0x8163: '…' // U+2026 HORIZONTAL ELLIPSIS
	0x8164: '‥' // U+2025 TWO DOT LEADER
	0x8165: '‘' // U+2018 LEFT SINGLE QUOTATION MARK
	0x8166: '’' // U+2019 RIGHT SINGLE QUOTATION MARK
	0x8167: '“' // U+201C LEFT DOUBLE QUOTATION MARK
	0x8168: '”' // U+201D RIGHT DOUBLE QUOTATION MARK
	0x8169: '（' // U+FF08 FULLWIDTH LEFT PARENTHESIS
	0x816A: '）' // U+FF09 FULLWIDTH RIGHT PARENTHESIS
	0x816B: '〔' // U+3014 LEFT TORTOISE SHELL BRACKET
	0x816C: '〕' // U+3015 RIGHT TORTOISE SHELL BRACKET
	0x816D: '［' // U+FF3B FULLWIDTH LEFT SQUARE BRACKET
	0x816E: '］' // U+FF3D FULLWIDTH RIGHT SQUARE BRACKET
	0x816F: '｛' // U+FF5B FULLWIDTH LEFT CURLY BRACKET
	0x8170: '｝' // U+FF5D FULLWIDTH RIGHT CURLY BRACKET
	0x8171: '〈' // U+3008 LEFT ANGLE BRACKET
	0x8172: '〉' // U+3009 RIGHT ANGLE BRACKET
	0x8173: '《' // U+300A LEFT DOUBLE ANGLE BRACKET
	0x8174: '》' // U+300B RIGHT DOUBLE ANGLE BRACKET
	0x8175: '「' // U+300C LEFT CORNER BRACKET
	0x8176: '」' // U+300D RIGHT CORNER BRACKET
	0x8177: '『' // U+300E LEFT WHITE CORNER BRACKET
	0x8178: '』' // U+300F RIGHT WHITE CORNER BRACKET
	0x8179: '【' // U+3010 LEFT BLACK LENTICULAR BRACKET
	0x817A: '】' // U+3011 RIGHT BLACK LENTICULAR BRACKET
	0x817B: '＋' // U+FF0B FULLWIDTH PLUS SIGN
	0x817C: '−' // U+2212 MINUS SIGN
	0x817D: '±' // U+00B1 PLUS-MINUS SIGN
	0x817E: '×' // U+00D7 MULTIPLICATION SIGN
	0x8180: '÷' // U+00F7 DIVISION SIGN
	0x8181: '＝' // U+FF1D FULLWIDTH EQUALS SIGN
	0x8182: '≠' // U+2260 NOT EQUAL TO
	0x8183: '＜' // U+FF1C FULLWIDTH LESS-THAN SIGN
	0x8184: '＞' // U+FF1E FULLWIDTH GREATER-THAN SIGN
	0x8185: '≦' // U+2266 LESS-THAN OVER EQUAL TO
	0x8186: '≧' // U+2267 GREATER-THAN OVER EQUAL TO
	0x8187: '∞' // U+221E INFINITY
	0x8188: '∴' // U+2234 THEREFORE
	0x8189: '♂' // U+2642 MALE SIGN
	0x818A: '♀' // U+2640 FEMALE SIGN
	0x818B: '°' // U+00B0 DEGREE SIGN
	0x818C: '′' // U+2032 PRIME
	0x818D: '″' // U+2033 DOUBLE PRIME
	0x818E: '℃' // U+2103 DEGREE CELSIUS
	0x818F: '￥' // U+FFE5 FULLWIDTH YEN SIGN
	0x8190: '＄' // U+FF04 FULLWIDTH DOLLAR SIGN
	0x8191: '¢' // U+00A2 CENT SIGN
	0x8192: '£' // U+00A3 POUND SIGN
	0x8193: '％' // U+FF05 FULLWIDTH PERCENT SIGN
	0x8194: '＃' // U+FF03 FULLWIDTH NUMBER SIGN
	0x8195: '＆' // U+FF06 FULLWIDTH AMPERSAND
	0x8196: '＊' // U+FF0A FULLWIDTH ASTERISK
	0x8197: '＠' // U+FF20 FULLWIDTH COMMERCIAL AT
	0x8198: '§' // U+00A7 SECTION SIGN
	0x8199: '☆' // U+2606 WHITE STAR
	0x819A: '★' // U+2605 BLACK STAR
	0x819B: '○' // U+25CB WHITE CIRCLE
	0x819C: '●' // U+25CF BLACK CIRCLE
	0x819D: '◎' // U+25CE BULLSEYE
	0x819E: '◇' // U+25C7 WHITE DIAMOND
	0x819F: '◆' // U+25C6 BLACK DIAMOND
	0x81A0: '□' // U+25A1 WHITE SQUARE
	0x81A1: '■' // U+25A0 BLACK SQUARE
	0x81A2: '△' // U+25B3 WHITE UP-POINTING TRIANGLE
	0x81A3: '▲' // U+25B2 BLACK UP-POINTING TRIANGLE
	0x81A4: '▽' // U+25BD WHITE DOWN-POINTING TRIANGLE
	0x81A5: '▼' // U+25BC BLACK DOWN-POINTING TRIANGLE
	0x81A6: '※' // U+203B REFERENCE MARK
	0x81A7: '〒' // U+3012 POSTAL MARK
	0x81A8: '→' // U+2192 RIGHTWARDS ARROW
	0x81A9: '←' // U+2190 LEFTWARDS ARROW
	0x81AA: '↑' // U+2191 UPWARDS ARROW
	0x81AB: '↓' // U+2193 DOWNWARDS ARROW
	0x81AC: '〓' // U+3013 GETA MARK
	0x81AD: '＇' // U+FF07 FULLWIDTH APOSTROPHE
	0x81AE: '＂' // U+FF02 FULLWIDTH QUOTATION MARK
	0x81AF: '－' // U+FF0D FULLWIDTH HYPHEN-MINUS
	0x81B0: '~' // U+007E TILDE
	0x81B1: '〳' // U+3033 VERTICAL KANA REPEAT MARK UPPER HALF
	0x81B2: '〴' // U+3034 VERTICAL KANA REPEAT WITH VOICED SOUND MARK UPPER HALF
	0x81B3: '〵' // U+3035 VERTICAL KANA REPEAT MARK LOWER HALF
	0x81B4: '〻' // U+303B VERTICAL IDEOGRAPHIC ITERATION MARK
	0x81B5: '〼' // U+303C MASU MARK
	0x81B6: 'ヿ' // U+30FF KATAKANA DIGRAPH KOTO
	0x81B7: 'ゟ' // U+309F HIRAGANA DIGRAPH YORI
	0x81B8: '∈' // U+2208 ELEMENT OF
	0x81B9: '∋' // U+220B CONTAINS AS MEMBER
	0x81BA: '⊆' // U+2286 SUBSET OF OR EQUAL TO
	0x81BB: '⊇' // U+2287 SUPERSET OF OR EQUAL TO
	0x81BC: '⊂' // U+2282 SUBSET OF
	0x81BD: '⊃' // U+2283 SUPERSET OF
	0x81BE: '∪' // U+222A UNION
	0x81BF: '∩' // U+2229 INTERSECTION
	0x81C0: '⊄' // U+2284 NOT A SUBSET OF
	0x81C1: '⊅' // U+2285 NOT A SUPERSET OF
	0x81C2: '⊊' // U+228A SUBSET OF WITH NOT EQUAL TO
	0x81C3: '⊋' // U+228B SUPERSET OF WITH NOT EQUAL TO
	0x81C4: '∉' // U+2209 NOT AN ELEMENT OF
	0x81C5: '∅' // U+2205 EMPTY SET
	0x81C6: '⌅' // U+2305 PROJECTIVE
	0x81C7: '⌆' // U+2306 PERSPECTIVE
	0x81C8: '∧' // U+2227 LOGICAL AND
	0x81C9: '∨' // U+2228 LOGICAL OR
	0x81CA: '¬' // U+00AC NOT SIGN
	0x81CB: '⇒' // U+21D2 RIGHTWARDS DOUBLE ARROW
	0x81CC: '⇔' // U+21D4 LEFT RIGHT DOUBLE ARROW
	0x81CD: '∀' // U+2200 FOR ALL
	0x81CE: '∃' // U+2203 THERE EXISTS
	0x81CF: '⊕' // U+2295 CIRCLED PLUS
	0x81D0: '⊖' // U+2296 CIRCLED MINUS
	0x81D1: '⊗' // U+2297 CIRCLED TIMES
	0x81D2: '∥' // U+2225 PARALLEL TO
	0x81D3: '∦' // U+2226 NOT PARALLEL TO
	0x81D4: '｟' // U+FF5F FULLWIDTH LEFT WHITE PARENTHESIS
	0x81D5: '｠' // U+FF60 FULLWIDTH RIGHT WHITE PARENTHESIS
	0x81D6: '〘' // U+3018 LEFT WHITE TORTOISE SHELL BRACKET
	0x81D7: '〙' // U+3019 RIGHT WHITE TORTOISE SHELL BRACKET
	0x81D8: '〖' // U+3016 LEFT WHITE LENTICULAR BRACKET
	0x81D9: '〗' // U+3017 RIGHT WHITE LENTICULAR BRACKET
	0x81DA: '∠' // U+2220 ANGLE
	0x81DB: '⊥' // U+22A5 UP TACK
	0x81DC: '⌒' // U+2312 ARC
	0x81DD: '∂' // U+2202 PARTIAL DIFFERENTIAL
	0x81DE: '∇' // U+2207 NABLA
	0x81DF: '≡' // U+2261 IDENTICAL TO
	0x81E0: '≒' // U+2252 APPROXIMATELY EQUAL TO OR THE IMAGE OF
	0x81E1: '≪' // U+226A MUCH LESS-THAN
	0x81E2: '≫' // U+226B MUCH GREATER-THAN
	0x81E3: '√' // U+221A SQUARE ROOT
	0x81E4: '∽' // U+223D REVERSED TILDE
	0x81E5: '∝' // U+221D PROPORTIONAL TO
	0x81E6: '∵' // U+2235 BECAUSE
	0x81E7: '∫' // U+222B INTEGRAL
	0x81E8: '∬' // U+222C DOUBLE INTEGRAL
	0x81E9: '≢' // U+2262 NOT IDENTICAL TO
	0x81EA: '≃' // U+2243 ASYMPTOTICALLY EQUAL TO
	0x81EB: '≅' // U+2245 APPROXIMATELY EQUAL TO
	0x81EC: '≈' // U+2248 ALMOST EQUAL TO
	0x81ED: '≶' // U+2276 LESS-THAN OR GREATER-THAN
	0x81EE: '≷' // U+2277 GREATER-THAN OR LESS-THAN
	0x81EF: '↔' // U+2194 LEFT RIGHT ARROW
	0x81F0: 'Å' // U+212B ANGSTROM SIGN
	0x81F1: '‰' // U+2030 PER MILLE SIGN
	0x81F2: '♯' // U+266F MUSIC SHARP SIGN
	0x81F3: '♭' // U+266D MUSIC FLAT SIGN
	0x81F4: '♪' // U+266A EIGHTH NOTE
	0x81F5: '†' // U+2020 DAGGER
	0x81F6: '‡' // U+2021 DOUBLE DAGGER
	0x81F7: '¶' // U+00B6 PILCROW SIGN
	0x81F8: '♮' // U+266E MUSIC NATURAL SIGN
	0x81F9: '♫' // U+266B BEAMED EIGHTH NOTES
	0x81FA: '♬' // U+266C BEAMED SIXTEENTH NOTES
	0x81FB: '♩' // U+2669 QUARTER NOTE
	0x81FC: '◯' // U+25EF LARGE CIRCLE
	0x8240: '▷' // U+25B7 WHITE RIGHT-POINTING TRIANGLE
	0x8241: '▶' // U+25B6 BLACK RIGHT-POINTING TRIANGLE
	0x8242: '◁' // U+25C1 WHITE LEFT-POINTING TRIANGLE
	0x8243: '◀' // U+25C0 BLACK LEFT-POINTING TRIANGLE
	0x8244: '↗' // U+2197 NORTH EAST ARROW
	0x8245: '↘' // U+2198 SOUTH EAST ARROW
	0x8246: '↖' // U+2196 NORTH WEST ARROW
	0x8247: '↙' // U+2199 SOUTH WEST ARROW
	0x8248: '⇄' // U+21C4 RIGHTWARDS ARROW OVER LEFTWARDS ARROW
	0x8249: '⇨' // U+21E8 RIGHTWARDS WHITE ARROW
	0x824A: '⇦' // U+21E6 LEFTWARDS WHITE ARROW
	0x824B: '⇧' // U+21E7 UPWARDS WHITE ARROW
	0x824C: '⇩' // U+21E9 DOWNWARDS WHITE ARROW
	0x824D: '⤴' // U+2934 ARROW POINTING RIGHTWARDS THEN CURVING UPWARDS
	0x824E: '⤵' // U+2935 ARROW POINTING RIGHTWARDS THEN CURVING DOWNWARDS
	0x824F: '０' // U+FF10 FULLWIDTH DIGIT ZERO
	0x8250: '１' // U+FF11 FULLWIDTH DIGIT ONE
	0x8251: '２' // U+FF12 FULLWIDTH DIGIT TWO
	0x8252: '３' // U+FF13 FULLWIDTH DIGIT THREE
	0x8253: '４' // U+FF14 FULLWIDTH DIGIT FOUR
	0x8254: '５' // U+FF15 FULLWIDTH DIGIT FIVE
	0x8255: '６' // U+FF16 FULLWIDTH DIGIT SIX
	0x8256: '７' // U+FF17 FULLWIDTH DIGIT SEVEN
	0x8257: '８' // U+FF18 FULLWIDTH DIGIT EIGHT
	0x8258: '９' // U+FF19 FULLWIDTH DIGIT NINE
	0x8259: '⦿' // U+29BF CIRCLED BULLET
	0x825A: '◉' // U+25C9 FISHEYE
	0x825B: '〽' // U+303D PART ALTERNATION MARK
	0x825C: '﹆' // U+FE46 WHITE SESAME DOT
	0x825D: '﹅' // U+FE45 SESAME DOT
	0x825E: '◦' // U+25E6 WHITE BULLET
	0x825F: '•' // U+2022 BULLET
	0x8260: 'Ａ' // U+FF21 FULLWIDTH LATIN CAPITAL LETTER A
	0x8261: 'Ｂ' // U+FF22 FULLWIDTH LATIN CAPITAL LETTER B
	0x8262: 'Ｃ' // U+FF23 FULLWIDTH LATIN CAPITAL LETTER C
	0x8263: 'Ｄ' // U+FF24 FULLWIDTH LATIN CAPITAL LETTER D
	0x8264: 'Ｅ' // U+FF25 FULLWIDTH LATIN CAPITAL LETTER E
	0x8265: 'Ｆ' // U+FF26 FULLWIDTH LATIN CAPITAL LETTER F
	0x8266: 'Ｇ' // U+FF27 FULLWIDTH LATIN CAPITAL LETTER G
	0x8267: 'Ｈ' // U+FF28 FULLWIDTH LATIN CAPITAL LETTER H
	0x8268: 'Ｉ' // U+FF29 FULLWIDTH LATIN CAPITAL LETTER I
	0x8269: 'Ｊ' // U+FF2A FULLWIDTH LATIN CAPITAL LETTER J
	0x826A: 'Ｋ' // U+FF2B FULLWIDTH LATIN CAPITAL LETTER K
	0x826B: 'Ｌ' // U+FF2C FULLWIDTH LATIN CAPITAL LETTER L
	0x826C: 'Ｍ' // U+FF2D FULLWIDTH LATIN CAPITAL LETTER M
	0x826D: 'Ｎ' // U+FF2E FULLWIDTH LATIN CAPITAL LETTER N
	0x826E: 'Ｏ' // U+FF2F FULLWIDTH LATIN CAPITAL LETTER O
	0x826F: 'Ｐ' // U+FF30 FULLWIDTH LATIN CAPITAL LETTER P
	0x8270: 'Ｑ' // U+FF31 FULLWIDTH LATIN CAPITAL LETTER Q
	0x8271: 'Ｒ' // U+FF32 FULLWIDTH LATIN CAPITAL LETTER R
	0x8272: 'Ｓ' // U+FF33 FULLWIDTH LATIN CAPITAL LETTER S
	0x8273: 'Ｔ' // U+FF34 FULLWIDTH LATIN CAPITAL LETTER T
	0x8274: 'Ｕ' // U+FF35 FULLWIDTH LATIN CAPITAL LETTER U
	0x8275: 'Ｖ' // U+FF36 FULLWIDTH LATIN CAPITAL LETTER V
	0x8276: 'Ｗ' // U+FF37 FULLWIDTH LATIN CAPITAL LETTER W
	0x8277: 'Ｘ' // U+FF38 FULLWIDTH LATIN CAPITAL LETTER X
	0x8278: 'Ｙ' // U+FF39 FULLWIDTH LATIN CAPITAL LETTER Y
	0x8279: 'Ｚ' // U+FF3A FULLWIDTH LATIN CAPITAL LETTER Z
	0x827A: '∓' // U+2213 MINUS-OR-PLUS SIGN
	0x827B: 'ℵ' // U+2135 ALEF SYMBOL
	0x827C: 'ℏ' // U+210F PLANCK CONSTANT OVER TWO PI
	0x827D: '㏋' // U+33CB SQUARE HP
	0x827E: 'ℓ' // U+2113 SCRIPT SMALL L
	0x8280: '℧' // U+2127 INVERTED OHM SIGN
	0x8281: 'ａ' // U+FF41 FULLWIDTH LATIN SMALL LETTER A
	0x8282: 'ｂ' // U+FF42 FULLWIDTH LATIN SMALL LETTER B
	0x8283: 'ｃ' // U+FF43 FULLWIDTH LATIN SMALL LETTER C
	0x8284: 'ｄ' // U+FF44 FULLWIDTH LATIN SMALL LETTER D
	0x8285: 'ｅ' // U+FF45 FULLWIDTH LATIN SMALL LETTER E
	0x8286: 'ｆ' // U+FF46 FULLWIDTH LATIN SMALL LETTER F
	0x8287: 'ｇ' // U+FF47 FULLWIDTH LATIN SMALL LETTER G
	0x8288: 'ｈ' // U+FF48 FULLWIDTH LATIN SMALL LETTER H
	0x8289: 'ｉ' // U+FF49 FULLWIDTH LATIN SMALL LETTER I
	0x828A: 'ｊ' // U+FF4A FULLWIDTH LATIN SMALL LETTER J
	0x828B: 'ｋ' // U+FF4B FULLWIDTH LATIN SMALL LETTER K
	0x828C: 'ｌ' // U+FF4C FULLWIDTH LATIN SMALL LETTER L
	0x828D: 'ｍ' // U+FF4D FULLWIDTH LATIN SMALL LETTER M
	0x828E: 'ｎ' // U+FF4E FULLWIDTH LATIN SMALL LETTER N
	0x828F: 'ｏ' // U+FF4F FULLWIDTH LATIN SMALL LETTER O
	0x8290: 'ｐ' // U+FF50 FULLWIDTH LATIN SMALL LETTER P
	0x8291: 'ｑ' // U+FF51 FULLWIDTH LATIN SMALL LETTER Q
	0x8292: 'ｒ' // U+FF52 FULLWIDTH LATIN SMALL LETTER R
	0x8293: 'ｓ' // U+FF53 FULLWIDTH LATIN SMALL LETTER S
	0x8294: 'ｔ' // U+FF54 FULLWIDTH LATIN SMALL LETTER T
	0x8295: 'ｕ' // U+FF55 FULLWIDTH LATIN SMALL LETTER U
	0x8296: 'ｖ' // U+FF56 FULLWIDTH LATIN SMALL LETTER V
	0x8297: 'ｗ' // U+FF57 FULLWIDTH LATIN SMALL LETTER W
	0x8298: 'ｘ' // U+FF58 FULLWIDTH LATIN SMALL LETTER X
	0x8299: 'ｙ' // U+FF59 FULLWIDTH LATIN SMALL LETTER Y
	0x829A: 'ｚ' // U+FF5A FULLWIDTH LATIN SMALL LETTER Z
	0x829B: '゠' // U+30A0 KATAKANA-HIRAGANA DOUBLE HYPHEN
	0x829C: '–' // U+2013 EN DASH
	0x829D: '⧺' // U+29FA DOUBLE PLUS
	0x829E: '⧻' // U+29FB TRIPLE PLUS
	0x829F: 'ぁ' // U+3041 HIRAGANA LETTER SMALL A
	0x82A0: 'あ' // U+3042 HIRAGANA LETTER A
	0x82A1: 'ぃ' // U+3043 HIRAGANA LETTER SMALL I
	0x82A2: 'い' // U+3044 HIRAGANA LETTER I
	0x82A3: 'ぅ' // U+3045 HIRAGANA LETTER SMALL U
	0x82A4: 'う' // U+3046 HIRAGANA LETTER U
	0x82A5: 'ぇ' // U+3047 HIRAGANA LETTER SMALL E
	0x82A6: 'え' // U+3048 HIRAGANA LETTER E
	0x82A7: 'ぉ' // U+3049 HIRAGANA LETTER SMALL O
	0x82A8: 'お' // U+304A HIRAGANA LETTER O
	0x82A9: 'か' // U+304B HIRAGANA LETTER KA
	0x82AA: 'が' // U+304C HIRAGANA LETTER GA
	0x82AB: 'き' // U+304D HIRAGANA LETTER KI
	0x82AC: 'ぎ' // U+304E HIRAGANA LETTER GI
	0x82AD: 'く' // U+304F HIRAGANA LETTER KU
	0x82AE: 'ぐ' // U+3050 HIRAGANA LETTER GU
	0x82AF: 'け' // U+3051 HIRAGANA LETTER KE
	0x82B0: 'げ' // U+3052 HIRAGANA LETTER GE
	0x82B1: 'こ' // U+3053 HIRAGANA LETTER KO
	0x82B2: 'ご' // U+3054 HIRAGANA LETTER GO
	0x82B3: 'さ' // U+3055 HIRAGANA LETTER SA
	0x82B4: 'ざ' // U+3056 HIRAGANA LETTER ZA
	0x82B5: 'し' // U+3057 HIRAGANA LETTER SI
	0x82B6: 'じ' // U+3058 HIRAGANA LETTER ZI
	0x82B7: 'す' // U+3059 HIRAGANA LETTER SU
	0x82B8: 'ず' // U+305A HIRAGANA LETTER ZU
	0x82B9: 'せ' // U+305B HIRAGANA LETTER SE
	0x82BA: 'ぜ' // U+305C HIRAGANA LETTER ZE
	0x82BB: 'そ' // U+305D HIRAGANA LETTER SO
	0x82BC: 'ぞ' // U+305E HIRAGANA LETTER ZO
	0x82BD: 'た' // U+305F HIRAGANA LETTER TA
	0x82BE: 'だ' // U+3060 HIRAGANA LETTER DA
	0x82BF: 'ち' // U+3061 HIRAGANA LETTER TI
	0x82C0: 'ぢ' // U+3062 HIRAGANA LETTER DI
	0x82C1: 'っ' // U+3063 HIRAGANA LETTER SMALL TU
	0x82C2: 'つ' // U+3064 HIRAGANA LETTER TU
	0x82C3: 'づ' // U+3065 HIRAGANA LETTER DU
	0x82C4: 'て' // U+3066 HIRAGANA LETTER TE
	0x82C5: 'で' // U+3067 HIRAGANA LETTER DE
	0x82C6: 'と' // U+3068 HIRAGANA LETTER TO
	0x82C7: 'ど' // U+3069 HIRAGANA LETTER DO
	0x82C8: 'な' // U+306A HIRAGANA LETTER NA
	0x82C9: 'に' // U+306B HIRAGANA LETTER NI
	0x82CA: 'ぬ' // U+306C HIRAGANA LETTER NU
	0x82CB: 'ね' // U+306D HIRAGANA LETTER NE
	0x82CC: 'の' // U+306E HIRAGANA LETTER NO
	0x82CD: 'は' // U+306F HIRAGANA LETTER HA
	0x82CE: 'ば' // U+3070 HIRAGANA LETTER BA
	0x82CF: 'ぱ' // U+3071 HIRAGANA LETTER PA
	0x82D0: 'ひ' // U+3072 HIRAGANA LETTER HI
	0x82D1: 'び' // U+3073 HIRAGANA LETTER BI
	0x82D2: 'ぴ' // U+3074 HIRAGANA LETTER PI
	0x82D3: 'ふ' // U+3075 HIRAGANA LETTER HU
	0x82D4: 'ぶ' // U+3076 HIRAGANA LETTER BU
	0x82D5: 'ぷ' // U+3077 HIRAGANA LETTER PU
	0x82D6: 'へ' // U+3078 HIRAGANA LETTER HE
	0x82D7: 'べ' // U+3079 HIRAGANA LETTER BE
	0x82D8: 'ぺ' // U+307A HIRAGANA LETTER PE
	0x82D9: 'ほ' // U+307B HIRAGANA LETTER HO
	0x82DA: 'ぼ' // U+307C HIRAGANA LETTER BO
	0x82DB: 'ぽ' // U+307D HIRAGANA LETTER PO
	0x82DC: 'ま' // U+307E HIRAGANA LETTER MA
	0x82DD: 'み' // U+307F HIRAGANA LETTER MI
	0x82DE: 'む' // U+3080 HIRAGANA LETTER MU
	0x82DF: 'め' // U+3081 HIRAGANA LETTER ME
	0x82E0: 'も' // U+3082 HIRAGANA LETTER MO
	0x82E1: 'ゃ' // U+3083 HIRAGANA LETTER SMALL YA
	0x82E2: 'や' // U+3084 HIRAGANA LETTER YA
	0x82E3: 'ゅ' // U+3085 HIRAGANA LETTER SMALL YU
	0x82E4: 'ゆ' // U+3086 HIRAGANA LETTER YU
	0x82E5: 'ょ' // U+3087 HIRAGANA LETTER SMALL YO
	0x82E6: 'よ' // U+3088 HIRAGANA LETTER YO
	0x82E7: 'ら' // U+3089 HIRAGANA LETTER RA
	0x82E8: 'り' // U+308A HIRAGANA LETTER RI
	0x82E9: 'る' // U+308B HIRAGANA LETTER RU
	0x82EA: 'れ' // U+308C HIRAGANA LETTER RE
	0x82EB: 'ろ' // U+308D HIRAGANA LETTER RO
	0x82EC: 'ゎ' // U+308E HIRAGANA LETTER SMALL WA
	0x82ED: 'わ' // U+308F HIRAGANA LETTER WA
	0x82EE: 'ゐ' // U+3090 HIRAGANA LETTER WI
	0x82EF: 'ゑ' // U+3091 HIRAGANA LETTER WE
	0x82F0: 'を' // U+3092 HIRAGANA LETTER WO
	0x82F1: 'ん' // U+3093 HIRAGANA LETTER N
	0x82F2: 'ゔ' // U+3094 HIRAGANA LETTER VU
	0x82F3: 'ゕ' // U+3095 HIRAGANA LETTER SMALL KA
	0x82F4: 'ゖ' // U+3096 HIRAGANA LETTER SMALL KE
	0x82F5: 'か゚' // U+304B+309A
	0x82F6: 'き゚' // U+304D+309A
	0x82F7: 'く゚' // U+304F+309A
	0x82F8: 'け゚' // U+3051+309A
	0x82F9: 'こ゚' // U+3053+309A
	0x8340: 'ァ' // U+30A1 KATAKANA LETTER SMALL A
	0x8341: 'ア' // U+30A2 KATAKANA LETTER A
	0x8342: 'ィ' // U+30A3 KATAKANA LETTER SMALL I
	0x8343: 'イ' // U+30A4 KATAKANA LETTER I
	0x8344: 'ゥ' // U+30A5 KATAKANA LETTER SMALL U
	0x8345: 'ウ' // U+30A6 KATAKANA LETTER U
	0x8346: 'ェ' // U+30A7 KATAKANA LETTER SMALL E
	0x8347: 'エ' // U+30A8 KATAKANA LETTER E
	0x8348: 'ォ' // U+30A9 KATAKANA LETTER SMALL O
	0x8349: 'オ' // U+30AA KATAKANA LETTER O
	0x834A: 'カ' // U+30AB KATAKANA LETTER KA
	0x834B: 'ガ' // U+30AC KATAKANA LETTER GA
	0x834C: 'キ' // U+30AD KATAKANA LETTER KI
	0x834D: 'ギ' // U+30AE KATAKANA LETTER GI
	0x834E: 'ク' // U+30AF KATAKANA LETTER KU
	0x834F: 'グ' // U+30B0 KATAKANA LETTER GU
	0x8350: 'ケ' // U+30B1 KATAKANA LETTER KE
	0x8351: 'ゲ' // U+30B2 KATAKANA LETTER GE
	0x8352: 'コ' // U+30B3 KATAKANA LETTER KO
	0x8353: 'ゴ' // U+30B4 KATAKANA LETTER GO
	0x8354: 'サ' // U+30B5 KATAKANA LETTER SA
	0x8355: 'ザ' // U+30B6 KATAKANA LETTER ZA
	0x8356: 'シ' // U+30B7 KATAKANA LETTER SI
	0x8357: 'ジ' // U+30B8 KATAKANA LETTER ZI
	0x8358: 'ス' // U+30B9 KATAKANA LETTER SU
	0x8359: 'ズ' // U+30BA KATAKANA LETTER ZU
	0x835A: 'セ' // U+30BB KATAKANA LETTER SE
	0x835B: 'ゼ' // U+30BC KATAKANA LETTER ZE
	0x835C: 'ソ' // U+30BD KATAKANA LETTER SO
	0x835D: 'ゾ' // U+30BE KATAKANA LETTER ZO
	0x835E: 'タ' // U+30BF KATAKANA LETTER TA
	0x835F: 'ダ' // U+30C0 KATAKANA LETTER DA
	0x8360: 'チ' // U+30C1 KATAKANA LETTER TI
	0x8361: 'ヂ' // U+30C2 KATAKANA LETTER DI
	0x8362: 'ッ' // U+30C3 KATAKANA LETTER SMALL TU
	0x8363: 'ツ' // U+30C4 KATAKANA LETTER TU
	0x8364: 'ヅ' // U+30C5 KATAKANA LETTER DU
	0x8365: 'テ' // U+30C6 KATAKANA LETTER TE
	0x8366: 'デ' // U+30C7 KATAKANA LETTER DE
	0x8367: 'ト' // U+30C8 KATAKANA LETTER TO
	0x8368: 'ド' // U+30C9 KATAKANA LETTER DO
	0x8369: 'ナ' // U+30CA KATAKANA LETTER NA
	0x836A: 'ニ' // U+30CB KATAKANA LETTER NI
	0x836B: 'ヌ' // U+30CC KATAKANA LETTER NU
	0x836C: 'ネ' // U+30CD KATAKANA LETTER NE
	0x836D: 'ノ' // U+30CE KATAKANA LETTER NO
	0x836E: 'ハ' // U+30CF KATAKANA LETTER HA
	0x836F: 'バ' // U+30D0 KATAKANA LETTER BA
	0x8370: 'パ' // U+30D1 KATAKANA LETTER PA
	0x8371: 'ヒ' // U+30D2 KATAKANA LETTER HI
	0x8372: 'ビ' // U+30D3 KATAKANA LETTER BI
	0x8373: 'ピ' // U+30D4 KATAKANA LETTER PI
	0x8374: 'フ' // U+30D5 KATAKANA LETTER HU
	0x8375: 'ブ' // U+30D6 KATAKANA LETTER BU
	0x8376: 'プ' // U+30D7 KATAKANA LETTER PU
	0x8377: 'ヘ' // U+30D8 KATAKANA LETTER HE
	0x8378: 'ベ' // U+30D9 KATAKANA LETTER BE
	0x8379: 'ペ' // U+30DA KATAKANA LETTER PE
	0x837A: 'ホ' // U+30DB KATAKANA LETTER HO
	0x837B: 'ボ' // U+30DC KATAKANA LETTER BO
	0x837C: 'ポ' // U+30DD KATAKANA LETTER PO
	0x837D: 'マ' // U+30DE KATAKANA LETTER MA
	0x837E: 'ミ' // U+30DF KATAKANA LETTER MI
	0x8380: 'ム' // U+30E0 KATAKANA LETTER MU
	0x8381: 'メ' // U+30E1 KATAKANA LETTER ME
	0x8382: 'モ' // U+30E2 KATAKANA LETTER MO
	0x8383: 'ャ' // U+30E3 KATAKANA LETTER SMALL YA
	0x8384: 'ヤ' // U+30E4 KATAKANA LETTER YA
	0x8385: 'ュ' // U+30E5 KATAKANA LETTER SMALL YU
	0x8386: 'ユ' // U+30E6 KATAKANA LETTER YU
	0x8387: 'ョ' // U+30E7 KATAKANA LETTER SMALL YO
	0x8388: 'ヨ' // U+30E8 KATAKANA LETTER YO
	0x8389: 'ラ' // U+30E9 KATAKANA LETTER RA
	0x838A: 'リ' // U+30EA KATAKANA LETTER RI
	0x838B: 'ル' // U+30EB KATAKANA LETTER RU
	0x838C: 'レ' // U+30EC KATAKANA LETTER RE
	0x838D: 'ロ' // U+30ED KATAKANA LETTER RO
	0x838E: 'ヮ' // U+30EE KATAKANA LETTER SMALL WA
	0x838F: 'ワ' // U+30EF KATAKANA LETTER WA
	0x8390: 'ヰ' // U+30F0 KATAKANA LETTER WI
	0x8391: 'ヱ' // U+30F1 KATAKANA LETTER WE
	0x8392: 'ヲ' // U+30F2 KATAKANA LETTER WO
	0x8393: 'ン' // U+30F3 KATAKANA LETTER N
	0x8394: 'ヴ' // U+30F4 KATAKANA LETTER VU
	0x8395: 'ヵ' // U+30F5 KATAKANA LETTER SMALL KA
	0x8396: 'ヶ' // U+30F6 KATAKANA LETTER SMALL KE
	0x8397: 'カ゚' // U+30AB+309A
	0x8398: 'キ゚' // U+30AD+309A
	0x8399: 'ク゚' // U+30AF+309A
	0x839A: 'ケ゚' // U+30B1+309A
	0x839B: 'コ゚' // U+30B3+309A
	0x839C: 'セ゚' // U+30BB+309A
	0x839D: 'ツ゚' // U+30C4+309A
	0x839E: 'ト゚' // U+30C8+309A
	0x839F: 'Α' // U+0391 GREEK CAPITAL LETTER ALPHA
	0x83A0: 'Β' // U+0392 GREEK CAPITAL LETTER BETA
	0x83A1: 'Γ' // U+0393 GREEK CAPITAL LETTER GAMMA
	0x83A2: 'Δ' // U+0394 GREEK CAPITAL LETTER DELTA
	0x83A3: 'Ε' // U+0395 GREEK CAPITAL LETTER EPSILON
	0x83A4: 'Ζ' // U+0396 GREEK CAPITAL LETTER ZETA
	0x83A5: 'Η' // U+0397 GREEK CAPITAL LETTER ETA
	0x83A6: 'Θ' // U+0398 GREEK CAPITAL LETTER THETA
	0x83A7: 'Ι' // U+0399 GREEK CAPITAL LETTER IOTA
	0x83A8: 'Κ' // U+039A GREEK CAPITAL LETTER KAPPA
	0x83A9: 'Λ' // U+039B GREEK CAPITAL LETTER LAMDA
	0x83AA: 'Μ' // U+039C GREEK CAPITAL LETTER MU
	0x83AB: 'Ν' // U+039D GREEK CAPITAL LETTER NU
	0x83AC: 'Ξ' // U+039E GREEK CAPITAL LETTER XI
	0x83AD: 'Ο' // U+039F GREEK CAPITAL LETTER OMICRON
	0x83AE: 'Π' // U+03A0 GREEK CAPITAL LETTER PI
	0x83AF: 'Ρ' // U+03A1 GREEK CAPITAL LETTER RHO
	0x83B0: 'Σ' // U+03A3 GREEK CAPITAL LETTER SIGMA
	0x83B1: 'Τ' // U+03A4 GREEK CAPITAL LETTER TAU
	0x83B2: 'Υ' // U+03A5 GREEK CAPITAL LETTER UPSILON
	0x83B3: 'Φ' // U+03A6 GREEK CAPITAL LETTER PHI
	0x83B4: 'Χ' // U+03A7 GREEK CAPITAL LETTER CHI
	0x83B5: 'Ψ' // U+03A8 GREEK CAPITAL LETTER PSI
	0x83B6: 'Ω' // U+03A9 GREEK CAPITAL LETTER OMEGA
	0x83B7: '♤' // U+2664 WHITE SPADE SUIT
	0x83B8: '♠' // U+2660 BLACK SPADE SUIT
	0x83B9: '♢' // U+2662 WHITE DIAMOND SUIT
	0x83BA: '♦' // U+2666 BLACK DIAMOND SUIT
	0x83BB: '♡' // U+2661 WHITE HEART SUIT
	0x83BC: '♥' // U+2665 BLACK HEART SUIT
	0x83BD: '♧' // U+2667 WHITE CLUB SUIT
	0x83BE: '♣' // U+2663 BLACK CLUB SUIT
	0x83BF: 'α' // U+03B1 GREEK SMALL LETTER ALPHA
	0x83C0: 'β' // U+03B2 GREEK SMALL LETTER BETA
	0x83C1: 'γ' // U+03B3 GREEK SMALL LETTER GAMMA
	0x83C2: 'δ' // U+03B4 GREEK SMALL LETTER DELTA
	0x83C3: 'ε' // U+03B5 GREEK SMALL LETTER EPSILON
	0x83C4: 'ζ' // U+03B6 GREEK SMALL LETTER ZETA
	0x83C5: 'η' // U+03B7 GREEK SMALL LETTER ETA
	0x83C6: 'θ' // U+03B8 GREEK SMALL LETTER THETA
	0x83C7: 'ι' // U+03B9 GREEK SMALL LETTER IOTA
	0x83C8: 'κ' // U+03BA GREEK SMALL LETTER KAPPA
	0x83C9: 'λ' // U+03BB GREEK SMALL LETTER LAMDA
	0x83CA: 'μ' // U+03BC GREEK SMALL LETTER MU
	0x83CB: 'ν' // U+03BD GREEK SMALL LETTER NU
	0x83CC: 'ξ' // U+03BE GREEK SMALL LETTER XI
	0x83CD: 'ο' // U+03BF GREEK SMALL LETTER OMICRON
	0x83CE: 'π' // U+03C0 GREEK SMALL LETTER PI
	0x83CF: 'ρ' // U+03C1 GREEK SMALL LETTER RHO
	0x83D0: 'σ' // U+03C3 GREEK SMALL LETTER SIGMA
	0x83D1: 'τ' // U+03C4 GREEK SMALL LETTER TAU
	0x83D2: 'υ' // U+03C5 GREEK SMALL LETTER UPSILON
	0x83D3: 'φ' // U+03C6 GREEK SMALL LETTER PHI
	0x83D4: 'χ' // U+03C7 GREEK SMALL LETTER CHI
	0x83D5: 'ψ' // U+03C8 GREEK SMALL LETTER PSI
	0x83D6: 'ω' // U+03C9 GREEK SMALL LETTER OMEGA
	0x83D7: 'ς' // U+03C2 GREEK SMALL LETTER FINAL SIGMA
	0x83D8: '⓵' // U+24F5 DOUBLE CIRCLED DIGIT ONE
	0x83D9: '⓶' // U+24F6 DOUBLE CIRCLED DIGIT TWO
	0x83DA: '⓷' // U+24F7 DOUBLE CIRCLED DIGIT THREE
	0x83DB: '⓸' // U+24F8 DOUBLE CIRCLED DIGIT FOUR
	0x83DC: '⓹' // U+24F9 DOUBLE CIRCLED DIGIT FIVE
	0x83DD: '⓺' // U+24FA DOUBLE CIRCLED DIGIT SIX
	0x83DE: '⓻' // U+24FB DOUBLE CIRCLED DIGIT SEVEN
	0x83DF: '⓼' // U+24FC DOUBLE CIRCLED DIGIT EIGHT
	0x83E0: '⓽' // U+24FD DOUBLE CIRCLED DIGIT NINE
	0x83E1: '⓾' // U+24FE DOUBLE CIRCLED NUMBER TEN
	0x83E2: '☖' // U+2616 WHITE SHOGI PIECE
	0x83E3: '☗' // U+2617 BLACK SHOGI PIECE
	0x83E4: '〠' // U+3020 POSTAL MARK FACE
	0x83E5: '☎' // U+260E BLACK TELEPHONE
	0x83E6: '☀' // U+2600 BLACK SUN WITH RAYS
	0x83E7: '☁' // U+2601 CLOUD
	0x83E8: '☂' // U+2602 UMBRELLA
	0x83E9: '☃' // U+2603 SNOWMAN
	0x83EA: '♨' // U+2668 HOT SPRINGS
	0x83EB: '▱' // U+25B1 WHITE PARALLELOGRAM
	0x83EC: 'ㇰ' // U+31F0 KATAKANA LETTER SMALL KU
	0x83ED: 'ㇱ' // U+31F1 KATAKANA LETTER SMALL SI
	0x83EE: 'ㇲ' // U+31F2 KATAKANA LETTER SMALL SU
	0x83EF: 'ㇳ' // U+31F3 KATAKANA LETTER SMALL TO
	0x83F0: 'ㇴ' // U+31F4 KATAKANA LETTER SMALL NU
	0x83F1: 'ㇵ' // U+31F5 KATAKANA LETTER SMALL HA
	0x83F2: 'ㇶ' // U+31F6 KATAKANA LETTER SMALL HI
	0x83F3: 'ㇷ' // U+31F7 KATAKANA LETTER SMALL HU
	0x83F4: 'ㇸ' // U+31F8 KATAKANA LETTER SMALL HE
	0x83F5: 'ㇹ' // U+31F9 KATAKANA LETTER SMALL HO
	0x83F6: 'ㇷ゚' // U+31F7+309A
	0x83F7: 'ㇺ' // U+31FA KATAKANA LETTER SMALL MU
	0x83F8: 'ㇻ' // U+31FB KATAKANA LETTER SMALL RA
	0x83F9: 'ㇼ' // U+31FC KATAKANA LETTER SMALL RI
	0x83FA: 'ㇽ' // U+31FD KATAKANA LETTER SMALL RU
	0x83FB: 'ㇾ' // U+31FE KATAKANA LETTER SMALL RE
	0x83FC: 'ㇿ' // U+31FF KATAKANA LETTER SMALL RO
	0x8440: 'А' // U+0410 CYRILLIC CAPITAL LETTER A
	0x8441: 'Б' // U+0411 CYRILLIC CAPITAL LETTER BE
	0x8442: 'В' // U+0412 CYRILLIC CAPITAL LETTER VE
	0x8443: 'Г' // U+0413 CYRILLIC CAPITAL LETTER GHE
	0x8444: 'Д' // U+0414 CYRILLIC CAPITAL LETTER DE
	0x8445: 'Е' // U+0415 CYRILLIC CAPITAL LETTER IE
	0x8446: 'Ё' // U+0401 CYRILLIC CAPITAL LETTER IO
	0x8447: 'Ж' // U+0416 CYRILLIC CAPITAL LETTER ZHE
	0x8448: 'З' // U+0417 CYRILLIC CAPITAL LETTER ZE
	0x8449: 'И' // U+0418 CYRILLIC CAPITAL LETTER I
	0x844A: 'Й' // U+0419 CYRILLIC CAPITAL LETTER SHORT I
	0x844B: 'К' // U+041A CYRILLIC CAPITAL LETTER KA
	0x844C: 'Л' // U+041B CYRILLIC CAPITAL LETTER EL
	0x844D: 'М' // U+041C CYRILLIC CAPITAL LETTER EM
	0x844E: 'Н' // U+041D CYRILLIC CAPITAL LETTER EN
	0x844F: 'О' // U+041E CYRILLIC CAPITAL LETTER O
	0x8450: 'П' // U+041F CYRILLIC CAPITAL LETTER PE
	0x8451: 'Р' // U+0420 CYRILLIC CAPITAL LETTER ER
	0x8452: 'С' // U+0421 CYRILLIC CAPITAL LETTER ES
	0x8453: 'Т' // U+0422 CYRILLIC CAPITAL LETTER TE
	0x8454: 'У' // U+0423 CYRILLIC CAPITAL LETTER U
	0x8455: 'Ф' // U+0424 CYRILLIC CAPITAL LETTER EF
	0x8456: 'Х' // U+0425 CYRILLIC CAPITAL LETTER HA
	0x8457: 'Ц' // U+0426 CYRILLIC CAPITAL LETTER TSE
	0x8458: 'Ч' // U+0427 CYRILLIC CAPITAL LETTER CHE
	0x8459: 'Ш' // U+0428 CYRILLIC CAPITAL LETTER SHA
	0x845A: 'Щ' // U+0429 CYRILLIC CAPITAL LETTER SHCHA
	0x845B: 'Ъ' // U+042A CYRILLIC CAPITAL LETTER HARD SIGN
	0x845C: 'Ы' // U+042B CYRILLIC CAPITAL LETTER YERU
	0x845D: 'Ь' // U+042C CYRILLIC CAPITAL LETTER SOFT SIGN
	0x845E: 'Э' // U+042D CYRILLIC CAPITAL LETTER E
	0x845F: 'Ю' // U+042E CYRILLIC CAPITAL LETTER YU
	0x8460: 'Я' // U+042F CYRILLIC CAPITAL LETTER YA
	0x8461: '⎾' // U+23BE DENTISTRY SYMBOL LIGHT VERTICAL AND TOP RIGHT
	0x8462: '⎿' // U+23BF DENTISTRY SYMBOL LIGHT VERTICAL AND BOTTOM RIGHT
	0x8463: '⏀' // U+23C0 DENTISTRY SYMBOL LIGHT VERTICAL WITH CIRCLE
	0x8464: '⏁' // U+23C1 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL WITH CIRCLE
	0x8465: '⏂' // U+23C2 DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL WITH CIRCLE
	0x8466: '⏃' // U+23C3 DENTISTRY SYMBOL LIGHT VERTICAL WITH TRIANGLE
	0x8467: '⏄' // U+23C4 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL WITH TRIANGLE
	0x8468: '⏅' // U+23C5 DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL WITH TRIANGLE
	0x8469: '⏆' // U+23C6 DENTISTRY SYMBOL LIGHT VERTICAL AND WAVE
	0x846A: '⏇' // U+23C7 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL WITH WAVE
	0x846B: '⏈' // U+23C8 DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL WITH WAVE
	0x846C: '⏉' // U+23C9 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL
	0x846D: '⏊' // U+23CA DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL
	0x846E: '⏋' // U+23CB DENTISTRY SYMBOL LIGHT VERTICAL AND TOP LEFT
	0x846F: '⏌' // U+23CC DENTISTRY SYMBOL LIGHT VERTICAL AND BOTTOM LEFT
	0x8470: 'а' // U+0430 CYRILLIC SMALL LETTER A
	0x8471: 'б' // U+0431 CYRILLIC SMALL LETTER BE
	0x8472: 'в' // U+0432 CYRILLIC SMALL LETTER VE
	0x8473: 'г' // U+0433 CYRILLIC SMALL LETTER GHE
	0x8474: 'д' // U+0434 CYRILLIC SMALL LETTER DE
	0x8475: 'е' // U+0435 CYRILLIC SMALL LETTER IE
	0x8476: 'ё' // U+0451 CYRILLIC SMALL LETTER IO
	0x8477: 'ж' // U+0436 CYRILLIC SMALL LETTER ZHE
	0x8478: 'з' // U+0437 CYRILLIC SMALL LETTER ZE
	0x8479: 'и' // U+0438 CYRILLIC SMALL LETTER I
	0x847A: 'й' // U+0439 CYRILLIC SMALL LETTER SHORT I
	0x847B: 'к' // U+043A CYRILLIC SMALL LETTER KA
	0x847C: 'л' // U+043B CYRILLIC SMALL LETTER EL
	0x847D: 'м' // U+043C CYRILLIC SMALL LETTER EM
	0x847E: 'н' // U+043D CYRILLIC SMALL LETTER EN
	0x8480: 'о' // U+043E CYRILLIC SMALL LETTER O
	0x8481: 'п' // U+043F CYRILLIC SMALL LETTER PE
	0x8482: 'р' // U+0440 CYRILLIC SMALL LETTER ER
	0x8483: 'с' // U+0441 CYRILLIC SMALL LETTER ES
	0x8484: 'т' // U+0442 CYRILLIC SMALL LETTER TE
	0x8485: 'у' // U+0443 CYRILLIC SMALL LETTER U
	0x8486: 'ф' // U+0444 CYRILLIC SMALL LETTER EF
	0x8487: 'х' // U+0445 CYRILLIC SMALL LETTER HA
	0x8488: 'ц' // U+0446 CYRILLIC SMALL LETTER TSE
	0x8489: 'ч' // U+0447 CYRILLIC SMALL LETTER CHE
	0x848A: 'ш' // U+0448 CYRILLIC SMALL LETTER SHA
	0x848B: 'щ' // U+0449 CYRILLIC SMALL LETTER SHCHA
	0x848C: 'ъ' // U+044A CYRILLIC SMALL LETTER HARD SIGN
	0x848D: 'ы' // U+044B CYRILLIC SMALL LETTER YERU
	0x848E: 'ь' // U+044C CYRILLIC SMALL LETTER SOFT SIGN
	0x848F: 'э' // U+044D CYRILLIC SMALL LETTER E
	0x8490: 'ю' // U+044E CYRILLIC SMALL LETTER YU
	0x8491: 'я' // U+044F CYRILLIC SMALL LETTER YA
	0x8492: 'ヷ' // U+30F7 KATAKANA LETTER VA
	0x8493: 'ヸ' // U+30F8 KATAKANA LETTER VI
	0x8494: 'ヹ' // U+30F9 KATAKANA LETTER VE
	0x8495: 'ヺ' // U+30FA KATAKANA LETTER VO
	0x8496: '⋚' // U+22DA LESS-THAN EQUAL TO OR GREATER-THAN
	0x8497: '⋛' // U+22DB GREATER-THAN EQUAL TO OR LESS-THAN
	0x8498: '⅓' // U+2153 VULGAR FRACTION ONE THIRD
	0x8499: '⅔' // U+2154 VULGAR FRACTION TWO THIRDS
	0x849A: '⅕' // U+2155 VULGAR FRACTION ONE FIFTH
	0x849B: '✓' // U+2713 CHECK MARK
	0x849C: '⌘' // U+2318 PLACE OF INTEREST SIGN
	0x849D: '␣' // U+2423 OPEN BOX
	0x849E: '⏎' // U+23CE RETURN SYMBOL
	0x849F: '─' // U+2500 BOX DRAWINGS LIGHT HORIZONTAL
	0x84A0: '│' // U+2502 BOX DRAWINGS LIGHT VERTICAL
	0x84A1: '┌' // U+250C BOX DRAWINGS LIGHT DOWN AND RIGHT
	0x84A2: '┐' // U+2510 BOX DRAWINGS LIGHT DOWN AND LEFT
	0x84A3: '┘' // U+2518 BOX DRAWINGS LIGHT UP AND LEFT
	0x84A4: '└' // U+2514 BOX DRAWINGS LIGHT UP AND RIGHT
	0x84A5: '├' // U+251C BOX DRAWINGS LIGHT VERTICAL AND RIGHT
	0x84A6: '┬' // U+252C BOX DRAWINGS LIGHT DOWN AND HORIZONTAL
	0x84A7: '┤' // U+2524 BOX DRAWINGS LIGHT VERTICAL AND LEFT
	0x84A8: '┴' // U+2534 BOX DRAWINGS LIGHT UP AND HORIZONTAL
	0x84A9: '┼' // U+253C BOX DRAWINGS LIGHT VERTICAL AND HORIZONTAL
	0x84AA: '━' // U+2501 BOX DRAWINGS HEAVY HORIZONTAL
	0x84AB: '┃' // U+2503 BOX DRAWINGS HEAVY VERTICAL
	0x84AC: '┏' // U+250F BOX DRAWINGS HEAVY DOWN AND RIGHT
	0x84AD: '┓' // U+2513 BOX DRAWINGS HEAVY DOWN AND LEFT
	0x84AE: '┛' // U+251B BOX DRAWINGS HEAVY UP AND LEFT
	0x84AF: '┗' // U+2517 BOX DRAWINGS HEAVY UP AND RIGHT
	0x84B0: '┣' // U+2523 BOX DRAWINGS HEAVY VERTICAL AND RIGHT
	0x84B1: '┳' // U+2533 BOX DRAWINGS HEAVY DOWN AND HORIZONTAL
	0x84B2: '┫' // U+252B BOX DRAWINGS HEAVY VERTICAL AND LEFT
	0x84B3: '┻' // U+253B BOX DRAWINGS HEAVY UP AND HORIZONTAL
	0x84B4: '╋' // U+254B BOX DRAWINGS HEAVY VERTICAL AND HORIZONTAL
	0x84B5: '┠' // U+2520 BOX DRAWINGS VERTICAL HEAVY AND RIGHT LIGHT
	0x84B6: '┯' // U+252F BOX DRAWINGS DOWN LIGHT AND HORIZONTAL HEAVY
	0x84B7: '┨' // U+2528 BOX DRAWINGS VERTICAL HEAVY AND LEFT LIGHT
	0x84B8: '┷' // U+2537 BOX DRAWINGS UP LIGHT AND HORIZONTAL HEAVY
	0x84B9: '┿' // U+253F BOX DRAWINGS VERTICAL LIGHT AND HORIZONTAL HEAVY
	0x84BA: '┝' // U+251D BOX DRAWINGS VERTICAL LIGHT AND RIGHT HEAVY
	0x84BB: '┰' // U+2530 BOX DRAWINGS DOWN HEAVY AND HORIZONTAL LIGHT
	0x84BC: '┥' // U+2525 BOX DRAWINGS VERTICAL LIGHT AND LEFT HEAVY
	0x84BD: '┸' // U+2538 BOX DRAWINGS UP HEAVY AND HORIZONTAL LIGHT
	0x84BE: '╂' // U+2542 BOX DRAWINGS VERTICAL HEAVY AND HORIZONTAL LIGHT
	0x84BF: '㉑' // U+3251 CIRCLED NUMBER TWENTY ONE
	0x84C0: '㉒' // U+3252 CIRCLED NUMBER TWENTY TWO
	0x84C1: '㉓' // U+3253 CIRCLED NUMBER TWENTY THREE
	0x84C2: '㉔' // U+3254 CIRCLED NUMBER TWENTY FOUR
	0x84C3: '㉕' // U+3255 CIRCLED NUMBER TWENTY FIVE
	0x84C4: '㉖' // U+3256 CIRCLED NUMBER TWENTY SIX
	0x84C5: '㉗' // U+3257 CIRCLED NUMBER TWENTY SEVEN
	0x84C6: '㉘' // U+3258 CIRCLED NUMBER TWENTY EIGHT
	0x84C7: '㉙' // U+3259 CIRCLED NUMBER TWENTY NINE
	0x84C8: '㉚' // U+325A CIRCLED NUMBER THIRTY
	0x84C9: '㉛' // U+325B CIRCLED NUMBER THIRTY ONE
	0x84CA: '㉜' // U+325C CIRCLED NUMBER THIRTY TWO
	0x84CB: '㉝' // U+325D CIRCLED NUMBER THIRTY THREE
	0x84CC: '㉞' // U+325E CIRCLED NUMBER THIRTY FOUR
	0x84CD: '㉟' // U+325F CIRCLED NUMBER THIRTY FIVE
	0x84CE: '㊱' // U+32B1 CIRCLED NUMBER THIRTY SIX
	0x84CF: '㊲' // U+32B2 CIRCLED NUMBER THIRTY SEVEN
	0x84D0: '㊳' // U+32B3 CIRCLED NUMBER THIRTY EIGHT
	0x84D1: '㊴' // U+32B4 CIRCLED NUMBER THIRTY NINE
	0x84D2: '㊵' // U+32B5 CIRCLED NUMBER FORTY
	0x84D3: '㊶' // U+32B6 CIRCLED NUMBER FORTY ONE
	0x84D4: '㊷' // U+32B7 CIRCLED NUMBER FORTY TWO
	0x84D5: '㊸' // U+32B8 CIRCLED NUMBER FORTY THREE
	0x84D6: '㊹' // U+32B9 CIRCLED NUMBER FORTY FOUR
	0x84D7: '㊺' // U+32BA CIRCLED NUMBER FORTY FIVE
	0x84D8: '㊻' // U+32BB CIRCLED NUMBER FORTY SIX
	0x84D9: '㊼' // U+32BC CIRCLED NUMBER FORTY SEVEN
	0x84DA: '㊽' // U+32BD CIRCLED NUMBER FORTY EIGHT
	0x84DB: '㊾' // U+32BE CIRCLED NUMBER FORTY NINE
	0x84DC: '㊿' // U+32BF CIRCLED NUMBER FIFTY
	0x84E5: '◐' // U+25D0 CIRCLE WITH LEFT HALF BLACK
	0x84E6: '◑' // U+25D1 CIRCLE WITH RIGHT HALF BLACK
	0x84E7: '◒' // U+25D2 CIRCLE WITH LOWER HALF BLACK
	0x84E8: '◓' // U+25D3 CIRCLE WITH UPPER HALF BLACK
	0x84E9: '‼' // U+203C DOUBLE EXCLAMATION MARK
	0x84EA: '⁇' // U+2047 DOUBLE QUESTION MARK
	0x84EB: '⁈' // U+2048 QUESTION EXCLAMATION MARK
	0x84EC: '⁉' // U+2049 EXCLAMATION QUESTION MARK
	0x84ED: 'Ǎ' // U+01CD LATIN CAPITAL LETTER A WITH CARON
	0x84EE: 'ǎ' // U+01CE LATIN SMALL LETTER A WITH CARON
	0x84EF: 'ǐ' // U+01D0 LATIN SMALL LETTER I WITH CARON
	0x84F0: 'Ḿ' // U+1E3E LATIN CAPITAL LETTER M WITH ACUTE
	0x84F1: 'ḿ' // U+1E3F LATIN SMALL LETTER M WITH ACUTE
	0x84F2: 'Ǹ' // U+01F8 LATIN CAPITAL LETTER N WITH GRAVE
	0x84F3: 'ǹ' // U+01F9 LATIN SMALL LETTER N WITH GRAVE
	0x84F4: 'Ǒ' // U+01D1 LATIN CAPITAL LETTER O WITH CARON
	0x84F5: 'ǒ' // U+01D2 LATIN SMALL LETTER O WITH CARON
	0x84F6: 'ǔ' // U+01D4 LATIN SMALL LETTER U WITH CARON
	0x84F7: 'ǖ' // U+01D6 LATIN SMALL LETTER U WITH DIAERESIS AND MACRON
	0x84F8: 'ǘ' // U+01D8 LATIN SMALL LETTER U WITH DIAERESIS AND ACUTE
	0x84F9: 'ǚ' // U+01DA LATIN SMALL LETTER U WITH DIAERESIS AND CARON
	0x84FA: 'ǜ' // U+01DC LATIN SMALL LETTER U WITH DIAERESIS AND GRAVE
	0x8540: '€' // U+20AC EURO SIGN
	0x8541: ' ' // U+00A0 NO-BREAK SPACE
	0x8542: '¡' // U+00A1 INVERTED EXCLAMATION MARK
	0x8543: '¤' // U+00A4 CURRENCY SIGN
	0x8544: '¦' // U+00A6 BROKEN BAR
	0x8545: '©' // U+00A9 COPYRIGHT SIGN
	0x8546: 'ª' // U+00AA FEMININE ORDINAL INDICATOR
	0x8547: '«' // U+00AB LEFT-POINTING DOUBLE ANGLE QUOTATION MARK
	0x8548: '­' // U+00AD SOFT HYPHEN
	0x8549: '®' // U+00AE REGISTERED SIGN
	0x854A: '¯' // U+00AF MACRON
	0x854B: '²' // U+00B2 SUPERSCRIPT TWO
	0x854C: '³' // U+00B3 SUPERSCRIPT THREE
	0x854D: '·' // U+00B7 MIDDLE DOT
	0x854E: '¸' // U+00B8 CEDILLA
	0x854F: '¹' // U+00B9 SUPERSCRIPT ONE
	0x8550: 'º' // U+00BA MASCULINE ORDINAL INDICATOR
	0x8551: '»' // U+00BB RIGHT-POINTING DOUBLE ANGLE QUOTATION MARK
	0x8552: '¼' // U+00BC VULGAR FRACTION ONE QUARTER
	0x8553: '½' // U+00BD VULGAR FRACTION ONE HALF
	0x8554: '¾' // U+00BE VULGAR FRACTION THREE QUARTERS
	0x8555: '¿' // U+00BF INVERTED QUESTION MARK
	0x8556: 'À' // U+00C0 LATIN CAPITAL LETTER A WITH GRAVE
	0x8557: 'Á' // U+00C1 LATIN CAPITAL LETTER A WITH ACUTE
	0x8558: 'Â' // U+00C2 LATIN CAPITAL LETTER A WITH CIRCUMFLEX
	0x8559: 'Ã' // U+00C3 LATIN CAPITAL LETTER A WITH TILDE
	0x855A: 'Ä' // U+00C4 LATIN CAPITAL LETTER A WITH DIAERESIS
	0x855B: 'Å' // U+00C5 LATIN CAPITAL LETTER A WITH RING ABOVE
	0x855C: 'Æ' // U+00C6 LATIN CAPITAL LETTER AE
	0x855D: 'Ç' // U+00C7 LATIN CAPITAL LETTER C WITH CEDILLA
	0x855E: 'È' // U+00C8 LATIN CAPITAL LETTER E WITH GRAVE
	0x855F: 'É' // U+00C9 LATIN CAPITAL LETTER E WITH ACUTE
	0x8560: 'Ê' // U+00CA LATIN CAPITAL LETTER E WITH CIRCUMFLEX
	0x8561: 'Ë' // U+00CB LATIN CAPITAL LETTER E WITH DIAERESIS
	0x8562: 'Ì' // U+00CC LATIN CAPITAL LETTER I WITH GRAVE
	0x8563: 'Í' // U+00CD LATIN CAPITAL LETTER I WITH ACUTE
	0x8564: 'Î' // U+00CE LATIN CAPITAL LETTER I WITH CIRCUMFLEX
	0x8565: 'Ï' // U+00CF LATIN CAPITAL LETTER I WITH DIAERESIS
	0x8566: 'Ð' // U+00D0 LATIN CAPITAL LETTER ETH
	0x8567: 'Ñ' // U+00D1 LATIN CAPITAL LETTER N WITH TILDE
	0x8568: 'Ò' // U+00D2 LATIN CAPITAL LETTER O WITH GRAVE
	0x8569: 'Ó' // U+00D3 LATIN CAPITAL LETTER O WITH ACUTE
	0x856A: 'Ô' // U+00D4 LATIN CAPITAL LETTER O WITH CIRCUMFLEX
	0x856B: 'Õ' // U+00D5 LATIN CAPITAL LETTER O WITH TILDE
	0x856C: 'Ö' // U+00D6 LATIN CAPITAL LETTER O WITH DIAERESIS
	0x856D: 'Ø' // U+00D8 LATIN CAPITAL LETTER O WITH STROKE
	0x856E: 'Ù' // U+00D9 LATIN CAPITAL LETTER U WITH GRAVE
	0x856F: 'Ú' // U+00DA LATIN CAPITAL LETTER U WITH ACUTE
	0x8570: 'Û' // U+00DB LATIN CAPITAL LETTER U WITH CIRCUMFLEX
	0x8571: 'Ü' // U+00DC LATIN CAPITAL LETTER U WITH DIAERESIS
	0x8572: 'Ý' // U+00DD LATIN CAPITAL LETTER Y WITH ACUTE
	0x8573: 'Þ' // U+00DE LATIN CAPITAL LETTER THORN
	0x8574: 'ß' // U+00DF LATIN SMALL LETTER SHARP S
	0x8575: 'à' // U+00E0 LATIN SMALL LETTER A WITH GRAVE
	0x8576: 'á' // U+00E1 LATIN SMALL LETTER A WITH ACUTE
	0x8577: 'â' // U+00E2 LATIN SMALL LETTER A WITH CIRCUMFLEX
	0x8578: 'ã' // U+00E3 LATIN SMALL LETTER A WITH TILDE
	0x8579: 'ä' // U+00E4 LATIN SMALL LETTER A WITH DIAERESIS
	0x857A: 'å' // U+00E5 LATIN SMALL LETTER A WITH RING ABOVE
	0x857B: 'æ' // U+00E6 LATIN SMALL LETTER AE
	0x857C: 'ç' // U+00E7 LATIN SMALL LETTER C WITH CEDILLA
	0x857D: 'è' // U+00E8 LATIN SMALL LETTER E WITH GRAVE
	0x857E: 'é' // U+00E9 LATIN SMALL LETTER E WITH ACUTE
	0x8580: 'ê' // U+00EA LATIN SMALL LETTER E WITH CIRCUMFLEX
	0x8581: 'ë' // U+00EB LATIN SMALL LETTER E WITH DIAERESIS
	0x8582: 'ì' // U+00EC LATIN SMALL LETTER I WITH GRAVE
	0x8583: 'í' // U+00ED LATIN SMALL LETTER I WITH ACUTE
	0x8584: 'î' // U+00EE LATIN SMALL LETTER I WITH CIRCUMFLEX
	0x8585: 'ï' // U+00EF LATIN SMALL LETTER I WITH DIAERESIS
	0x8586: 'ð' // U+00F0 LATIN SMALL LETTER ETH
	0x8587: 'ñ' // U+00F1 LATIN SMALL LETTER N WITH TILDE
	0x8588: 'ò' // U+00F2 LATIN SMALL LETTER O WITH GRAVE
	0x8589: 'ó' // U+00F3 LATIN SMALL LETTER O WITH ACUTE
	0x858A: 'ô' // U+00F4 LATIN SMALL LETTER O WITH CIRCUMFLEX
	0x858B: 'õ' // U+00F5 LATIN SMALL LETTER O WITH TILDE
	0x858C: 'ö' // U+00F6 LATIN SMALL LETTER O WITH DIAERESIS
	0x858D: 'ø' // U+00F8 LATIN SMALL LETTER O WITH STROKE
	0x858E: 'ù' // U+00F9 LATIN SMALL LETTER U WITH GRAVE
	0x858F: 'ú' // U+00FA LATIN SMALL LETTER U WITH ACUTE
	0x8590: 'û' // U+00FB LATIN SMALL LETTER U WITH CIRCUMFLEX
	0x8591: 'ü' // U+00FC LATIN SMALL LETTER U WITH DIAERESIS
	0x8592: 'ý' // U+00FD LATIN SMALL LETTER Y WITH ACUTE
	0x8593: 'þ' // U+00FE LATIN SMALL LETTER THORN
	0x8594: 'ÿ' // U+00FF LATIN SMALL LETTER Y WITH DIAERESIS
	0x8595: 'Ā' // U+0100 LATIN CAPITAL LETTER A WITH MACRON
	0x8596: 'Ī' // U+012A LATIN CAPITAL LETTER I WITH MACRON
	0x8597: 'Ū' // U+016A LATIN CAPITAL LETTER U WITH MACRON
	0x8598: 'Ē' // U+0112 LATIN CAPITAL LETTER E WITH MACRON
	0x8599: 'Ō' // U+014C LATIN CAPITAL LETTER O WITH MACRON
	0x859A: 'ā' // U+0101 LATIN SMALL LETTER A WITH MACRON
	0x859B: 'ī' // U+012B LATIN SMALL LETTER I WITH MACRON
	0x859C: 'ū' // U+016B LATIN SMALL LETTER U WITH MACRON
	0x859D: 'ē' // U+0113 LATIN SMALL LETTER E WITH MACRON
	0x859E: 'ō' // U+014D LATIN SMALL LETTER O WITH MACRON
	0x859F: 'Ą' // U+0104 LATIN CAPITAL LETTER A WITH OGONEK
	0x85A0: '˘' // U+02D8 BREVE
	0x85A1: 'Ł' // U+0141 LATIN CAPITAL LETTER L WITH STROKE
	0x85A2: 'Ľ' // U+013D LATIN CAPITAL LETTER L WITH CARON
	0x85A3: 'Ś' // U+015A LATIN CAPITAL LETTER S WITH ACUTE
	0x85A4: 'Š' // U+0160 LATIN CAPITAL LETTER S WITH CARON
	0x85A5: 'Ş' // U+015E LATIN CAPITAL LETTER S WITH CEDILLA
	0x85A6: 'Ť' // U+0164 LATIN CAPITAL LETTER T WITH CARON
	0x85A7: 'Ź' // U+0179 LATIN CAPITAL LETTER Z WITH ACUTE
	0x85A8: 'Ž' // U+017D LATIN CAPITAL LETTER Z WITH CARON
	0x85A9: 'Ż' // U+017B LATIN CAPITAL LETTER Z WITH DOT ABOVE
	0x85AA: 'ą' // U+0105 LATIN SMALL LETTER A WITH OGONEK
	0x85AB: '˛' // U+02DB OGONEK
	0x85AC: 'ł' // U+0142 LATIN SMALL LETTER L WITH STROKE
	0x85AD: 'ľ' // U+013E LATIN SMALL LETTER L WITH CARON
	0x85AE: 'ś' // U+015B LATIN SMALL LETTER S WITH ACUTE
	0x85AF: 'ˇ' // U+02C7 CARON
	0x85B0: 'š' // U+0161 LATIN SMALL LETTER S WITH CARON
	0x85B1: 'ş' // U+015F LATIN SMALL LETTER S WITH CEDILLA
	0x85B2: 'ť' // U+0165 LATIN SMALL LETTER T WITH CARON
	0x85B3: 'ź' // U+017A LATIN SMALL LETTER Z WITH ACUTE
	0x85B4: '˝' // U+02DD DOUBLE ACUTE ACCENT
	0x85B5: 'ž' // U+017E LATIN SMALL LETTER Z WITH CARON
	0x85B6: 'ż' // U+017C LATIN SMALL LETTER Z WITH DOT ABOVE
	0x85B7: 'Ŕ' // U+0154 LATIN CAPITAL LETTER R WITH ACUTE
	0x85B8: 'Ă' // U+0102 LATIN CAPITAL LETTER A WITH BREVE
	0x85B9: 'Ĺ' // U+0139 LATIN CAPITAL LETTER L WITH ACUTE
	0x85BA: 'Ć' // U+0106 LATIN CAPITAL LETTER C WITH ACUTE
	0x85BB: 'Č' // U+010C LATIN CAPITAL LETTER C WITH CARON
	0x85BC: 'Ę' // U+0118 LATIN CAPITAL LETTER E WITH OGONEK
	0x85BD: 'Ě' // U+011A LATIN CAPITAL LETTER E WITH CARON
	0x85BE: 'Ď' // U+010E LATIN CAPITAL LETTER D WITH CARON
	0x85BF: 'Ń' // U+0143 LATIN CAPITAL LETTER N WITH ACUTE
	0x85C0: 'Ň' // U+0147 LATIN CAPITAL LETTER N WITH CARON
	0x85C1: 'Ő' // U+0150 LATIN CAPITAL LETTER O WITH DOUBLE ACUTE
	0x85C2: 'Ř' // U+0158 LATIN CAPITAL LETTER R WITH CARON
	0x85C3: 'Ů' // U+016E LATIN CAPITAL LETTER U WITH RING ABOVE
	0x85C4: 'Ű' // U+0170 LATIN CAPITAL LETTER U WITH DOUBLE ACUTE
	0x85C5: 'Ţ' // U+0162 LATIN CAPITAL LETTER T WITH CEDILLA
	0x85C6: 'ŕ' // U+0155 LATIN SMALL LETTER R WITH ACUTE
	0x85C7: 'ă' // U+0103 LATIN SMALL LETTER A WITH BREVE
	0x85C8: 'ĺ' // U+013A LATIN SMALL LETTER L WITH ACUTE
	0x85C9: 'ć' // U+0107 LATIN SMALL LETTER C WITH ACUTE
	0x85CA: 'č' // U+010D LATIN SMALL LETTER C WITH CARON
	0x85CB: 'ę' // U+0119 LATIN SMALL LETTER E WITH OGONEK
	0x85CC: 'ě' // U+011B LATIN SMALL LETTER E WITH CARON
	0x85CD: 'ď' // U+010F LATIN SMALL LETTER D WITH CARON
	0x85CE: 'đ' // U+0111 LATIN SMALL LETTER D WITH STROKE
	0x85CF: 'ń' // U+0144 LATIN SMALL LETTER N WITH ACUTE
	0x85D0: 'ň' // U+0148 LATIN SMALL LETTER N WITH CARON
	0x85D1: 'ő' // U+0151 LATIN SMALL LETTER O WITH DOUBLE ACUTE
	0x85D2: 'ř' // U+0159 LATIN SMALL LETTER R WITH CARON
	0x85D3: 'ů' // U+016F LATIN SMALL LETTER U WITH RING ABOVE
	0x85D4: 'ű' // U+0171 LATIN SMALL LETTER U WITH DOUBLE ACUTE
	0x85D5: 'ţ' // U+0163 LATIN SMALL LETTER T WITH CEDILLA
	0x85D6: '˙' // U+02D9 DOT ABOVE
	0x85D7: 'Ĉ' // U+0108 LATIN CAPITAL LETTER C WITH CIRCUMFLEX
	0x85D8: 'Ĝ' // U+011C LATIN CAPITAL LETTER G WITH CIRCUMFLEX
	0x85D9: 'Ĥ' // U+0124 LATIN CAPITAL LETTER H WITH CIRCUMFLEX
	0x85DA: 'Ĵ' // U+0134 LATIN CAPITAL LETTER J WITH CIRCUMFLEX
	0x85DB: 'Ŝ' // U+015C LATIN CAPITAL LETTER S WITH CIRCUMFLEX
	0x85DC: 'Ŭ' // U+016C LATIN CAPITAL LETTER U WITH BREVE
	0x85DD: 'ĉ' // U+0109 LATIN SMALL LETTER C WITH CIRCUMFLEX
	0x85DE: 'ĝ' // U+011D LATIN SMALL LETTER G WITH CIRCUMFLEX
	0x85DF: 'ĥ' // U+0125 LATIN SMALL LETTER H WITH CIRCUMFLEX
	0x85E0: 'ĵ' // U+0135 LATIN SMALL LETTER J WITH CIRCUMFLEX
	0x85E1: 'ŝ' // U+015D LATIN SMALL LETTER S WITH CIRCUMFLEX
	0x85E2: 'ŭ' // U+016D LATIN SMALL LETTER U WITH BREVE
	0x85E3: 'ɱ' // U+0271 LATIN SMALL LETTER M WITH HOOK
	0x85E4: 'ʋ' // U+028B LATIN SMALL LETTER V WITH HOOK
	0x85E5: 'ɾ' // U+027E LATIN SMALL LETTER R WITH FISHHOOK
	0x85E6: 'ʃ' // U+0283 LATIN SMALL LETTER ESH
	0x85E7: 'ʒ' // U+0292 LATIN SMALL LETTER EZH
	0x85E8: 'ɬ' // U+026C LATIN SMALL LETTER L WITH BELT
	0x85E9: 'ɮ' // U+026E LATIN SMALL LETTER LEZH
	0x85EA: 'ɹ' // U+0279 LATIN SMALL LETTER TURNED R
	0x85EB: 'ʈ' // U+0288 LATIN SMALL LETTER T WITH RETROFLEX HOOK
	0x85EC: 'ɖ' // U+0256 LATIN SMALL LETTER D WITH TAIL
	0x85ED: 'ɳ' // U+0273 LATIN SMALL LETTER N WITH RETROFLEX HOOK
	0x85EE: 'ɽ' // U+027D LATIN SMALL LETTER R WITH TAIL
	0x85EF: 'ʂ' // U+0282 LATIN SMALL LETTER S WITH HOOK
	0x85F0: 'ʐ' // U+0290 LATIN SMALL LETTER Z WITH RETROFLEX HOOK
	0x85F1: 'ɻ' // U+027B LATIN SMALL LETTER TURNED R WITH HOOK
	0x85F2: 'ɭ' // U+026D LATIN SMALL LETTER L WITH RETROFLEX HOOK
	0x85F3: 'ɟ' // U+025F LATIN SMALL LETTER DOTLESS J WITH STROKE
	0x85F4: 'ɲ' // U+0272 LATIN SMALL LETTER N WITH LEFT HOOK
	0x85F5: 'ʝ' // U+029D LATIN SMALL LETTER J WITH CROSSED-TAIL
	0x85F6: 'ʎ' // U+028E LATIN SMALL LETTER TURNED Y
	0x85F7: 'ɡ' // U+0261 LATIN SMALL LETTER SCRIPT G
	0x85F8: 'ŋ' // U+014B LATIN SMALL LETTER ENG
	0x85F9: 'ɰ' // U+0270 LATIN SMALL LETTER TURNED M WITH LONG LEG
	0x85FA: 'ʁ' // U+0281 LATIN LETTER SMALL CAPITAL INVERTED R
	0x85FB: 'ħ' // U+0127 LATIN SMALL LETTER H WITH STROKE
	0x85FC: 'ʕ' // U+0295 LATIN LETTER PHARYNGEAL VOICED FRICATIVE
	0x8640: 'ʔ' // U+0294 LATIN LETTER GLOTTAL STOP
	0x8641: 'ɦ' // U+0266 LATIN SMALL LETTER H WITH HOOK
	0x8642: 'ʘ' // U+0298 LATIN LETTER BILABIAL CLICK
	0x8643: 'ǂ' // U+01C2 LATIN LETTER ALVEOLAR CLICK
	0x8644: 'ɓ' // U+0253 LATIN SMALL LETTER B WITH HOOK
	0x8645: 'ɗ' // U+0257 LATIN SMALL LETTER D WITH HOOK
	0x8646: 'ʄ' // U+0284 LATIN SMALL LETTER DOTLESS J WITH STROKE AND HOOK
	0x8647: 'ɠ' // U+0260 LATIN SMALL LETTER G WITH HOOK
	0x8648: 'Ɠ' // U+0193 LATIN CAPITAL LETTER G WITH HOOK
	0x8649: 'œ' // U+0153 LATIN SMALL LIGATURE OE
	0x864A: 'Œ' // U+0152 LATIN CAPITAL LIGATURE OE
	0x864B: 'ɨ' // U+0268 LATIN SMALL LETTER I WITH STROKE
	0x864C: 'ʉ' // U+0289 LATIN SMALL LETTER U BAR
	0x864D: 'ɘ' // U+0258 LATIN SMALL LETTER REVERSED E
	0x864E: 'ɵ' // U+0275 LATIN SMALL LETTER BARRED O
	0x864F: 'ə' // U+0259 LATIN SMALL LETTER SCHWA
	0x8650: 'ɜ' // U+025C LATIN SMALL LETTER REVERSED OPEN E
	0x8651: 'ɞ' // U+025E LATIN SMALL LETTER CLOSED REVERSED OPEN E
	0x8652: 'ɐ' // U+0250 LATIN SMALL LETTER TURNED A
	0x8653: 'ɯ' // U+026F LATIN SMALL LETTER TURNED M
	0x8654: 'ʊ' // U+028A LATIN SMALL LETTER UPSILON
	0x8655: 'ɤ' // U+0264 LATIN SMALL LETTER RAMS HORN
	0x8656: 'ʌ' // U+028C LATIN SMALL LETTER TURNED V
	0x8657: 'ɔ' // U+0254 LATIN SMALL LETTER OPEN O
	0x8658: 'ɑ' // U+0251 LATIN SMALL LETTER ALPHA
	0x8659: 'ɒ' // U+0252 LATIN SMALL LETTER TURNED ALPHA
	0x865A: 'ʍ' // U+028D LATIN SMALL LETTER TURNED W
	0x865B: 'ɥ' // U+0265 LATIN SMALL LETTER TURNED H
	0x865C: 'ʢ' // U+02A2 LATIN LETTER REVERSED GLOTTAL STOP WITH STROKE
	0x865D: 'ʡ' // U+02A1 LATIN LETTER GLOTTAL STOP WITH STROKE
	0x865E: 'ɕ' // U+0255 LATIN SMALL LETTER C WITH CURL
	0x865F: 'ʑ' // U+0291 LATIN SMALL LETTER Z WITH CURL
	0x8660: 'ɺ' // U+027A LATIN SMALL LETTER TURNED R WITH LONG LEG
	0x8661: 'ɧ' // U+0267 LATIN SMALL LETTER HENG WITH HOOK
	0x8662: 'ɚ' // U+025A LATIN SMALL LETTER SCHWA WITH HOOK
	0x8663: 'æ̀' // U+00E6+0300
	0x8664: 'ǽ' // U+01FD LATIN SMALL LETTER AE WITH ACUTE
	0x8665: 'ὰ' // U+1F70 GREEK SMALL LETTER ALPHA WITH VARIA
	0x8666: 'ά' // U+1F71 GREEK SMALL LETTER ALPHA WITH OXIA
	0x8667: 'ɔ̀' // U+0254+0300
	0x8668: 'ɔ́' // U+0254+0301
	0x8669: 'ʌ̀' // U+028C+0300
	0x866A: 'ʌ́' // U+028C+0301
	0x866B: 'ə̀' // U+0259+0300
	0x866C: 'ə́' // U+0259+0301
	0x866D: 'ɚ̀' // U+025A+0300
	0x866E: 'ɚ́' // U+025A+0301
	0x866F: 'ὲ' // U+1F72 GREEK SMALL LETTER EPSILON WITH VARIA
	0x8670: 'έ' // U+1F73 GREEK SMALL LETTER EPSILON WITH OXIA
	0x8671: '͡' // U+0361 COMBINING DOUBLE INVERTED BREVE
	0x8672: 'ˈ' // U+02C8 MODIFIER LETTER VERTICAL LINE
	0x8673: 'ˌ' // U+02CC MODIFIER LETTER LOW VERTICAL LINE
	0x8674: 'ː' // U+02D0 MODIFIER LETTER TRIANGULAR COLON
	0x8675: 'ˑ' // U+02D1 MODIFIER LETTER HALF TRIANGULAR COLON
	0x8676: '̆' // U+0306 COMBINING BREVE
	0x8677: '‿' // U+203F UNDERTIE
	0x8678: '̋' // U+030B COMBINING DOUBLE ACUTE ACCENT
	0x8679: '́' // U+0301 COMBINING ACUTE ACCENT
	0x867A: '̄' // U+0304 COMBINING MACRON
	0x867B: '̀' // U+0300 COMBINING GRAVE ACCENT
	0x867C: '̏' // U+030F COMBINING DOUBLE GRAVE ACCENT
	0x867D: '̌' // U+030C COMBINING CARON
	0x867E: '̂' // U+0302 COMBINING CIRCUMFLEX ACCENT
	0x8680: '˥' // U+02E5 MODIFIER LETTER EXTRA-HIGH TONE BAR
	0x8681: '˦' // U+02E6 MODIFIER LETTER HIGH TONE BAR
	0x8682: '˧' // U+02E7 MODIFIER LETTER MID TONE BAR
	0x8683: '˨' // U+02E8 MODIFIER LETTER LOW TONE BAR
	0x8684: '˩' // U+02E9 MODIFIER LETTER EXTRA-LOW TONE BAR
	0x8685: '˩˥' // U+02E9+02E5
	0x8686: '˥˩' // U+02E5+02E9
	0x8687: '̥' // U+0325 COMBINING RING BELOW
	0x8688: '̬' // U+032C COMBINING CARON BELOW
	0x8689: '̹' // U+0339 COMBINING RIGHT HALF RING BELOW
	0x868A: '̜' // U+031C COMBINING LEFT HALF RING BELOW
	0x868B: '̟' // U+031F COMBINING PLUS SIGN BELOW
	0x868C: '̠' // U+0320 COMBINING MINUS SIGN BELOW
	0x868D: '̈' // U+0308 COMBINING DIAERESIS
	0x868E: '̽' // U+033D COMBINING X ABOVE
	0x868F: '̩' // U+0329 COMBINING VERTICAL LINE BELOW
	0x8690: '̯' // U+032F COMBINING INVERTED BREVE BELOW
	0x8691: '˞' // U+02DE MODIFIER LETTER RHOTIC HOOK
	0x8692: '̤' // U+0324 COMBINING DIAERESIS BELOW
	0x8693: '̰' // U+0330 COMBINING TILDE BELOW
	0x8694: '̼' // U+033C COMBINING SEAGULL BELOW
	0x8695: '̴' // U+0334 COMBINING TILDE OVERLAY
	0x8696: '̝' // U+031D COMBINING UP TACK BELOW
	0x8697: '̞' // U+031E COMBINING DOWN TACK BELOW
	0x8698: '̘' // U+0318 COMBINING LEFT TACK BELOW
	0x8699: '̙' // U+0319 COMBINING RIGHT TACK BELOW
	0x869A: '̪' // U+032A COMBINING BRIDGE BELOW
	0x869B: '̺' // U+033A COMBINING INVERTED BRIDGE BELOW
	0x869C: '̻' // U+033B COMBINING SQUARE BELOW
	0x869D: '̃' // U+0303 COMBINING TILDE
	0x869E: '̚' // U+031A COMBINING LEFT ANGLE ABOVE
	0x869F: '❶' // U+2776 DINGBAT NEGATIVE CIRCLED DIGIT ONE
	0x86A0: '❷' // U+2777 DINGBAT NEGATIVE CIRCLED DIGIT TWO
	0x86A1: '❸' // U+2778 DINGBAT NEGATIVE CIRCLED DIGIT THREE
	0x86A2: '❹' // U+2779 DINGBAT NEGATIVE CIRCLED DIGIT FOUR
	0x86A3: '❺' // U+277A DINGBAT NEGATIVE CIRCLED DIGIT FIVE
	0x86A4: '❻' // U+277B DINGBAT NEGATIVE CIRCLED DIGIT SIX
	0x86A5: '❼' // U+277C DINGBAT NEGATIVE CIRCLED DIGIT SEVEN
	0x86A6: '❽' // U+277D DINGBAT NEGATIVE CIRCLED DIGIT EIGHT
	0x86A7: '❾' // U+277E DINGBAT NEGATIVE CIRCLED DIGIT NINE
	0x86A8: '❿' // U+277F DINGBAT NEGATIVE CIRCLED NUMBER TEN
	0x86A9: '⓫' // U+24EB NEGATIVE CIRCLED NUMBER ELEVEN
	0x86AA: '⓬' // U+24EC NEGATIVE CIRCLED NUMBER TWELVE
	0x86AB: '⓭' // U+24ED NEGATIVE CIRCLED NUMBER THIRTEEN
	0x86AC: '⓮' // U+24EE NEGATIVE CIRCLED NUMBER FOURTEEN
	0x86AD: '⓯' // U+24EF NEGATIVE CIRCLED NUMBER FIFTEEN
	0x86AE: '⓰' // U+24F0 NEGATIVE CIRCLED NUMBER SIXTEEN
	0x86AF: '⓱' // U+24F1 NEGATIVE CIRCLED NUMBER SEVENTEEN
	0x86B0: '⓲' // U+24F2 NEGATIVE CIRCLED NUMBER EIGHTEEN
	0x86B1: '⓳' // U+24F3 NEGATIVE CIRCLED NUMBER NINETEEN
	0x86B2: '⓴' // U+24F4 NEGATIVE CIRCLED NUMBER TWENTY
	0x86B3: 'ⅰ' // U+2170 SMALL ROMAN NUMERAL ONE
	0x86B4: 'ⅱ' // U+2171 SMALL ROMAN NUMERAL TWO
	0x86B5: 'ⅲ' // U+2172 SMALL ROMAN NUMERAL THREE
	0x86B6: 'ⅳ' // U+2173 SMALL ROMAN NUMERAL FOUR
	0x86B7: 'ⅴ' // U+2174 SMALL ROMAN NUMERAL FIVE
	0x86B8: 'ⅵ' // U+2175 SMALL ROMAN NUMERAL SIX
	0x86B9: 'ⅶ' // U+2176 SMALL ROMAN NUMERAL SEVEN
	0x86BA: 'ⅷ' // U+2177 SMALL ROMAN NUMERAL EIGHT
	0x86BB: 'ⅸ' // U+2178 SMALL ROMAN NUMERAL NINE
	0x86BC: 'ⅹ' // U+2179 SMALL ROMAN NUMERAL TEN
	0x86BD: 'ⅺ' // U+217A SMALL ROMAN NUMERAL ELEVEN
	0x86BE: 'ⅻ' // U+217B SMALL ROMAN NUMERAL TWELVE
	0x86BF: 'ⓐ' // U+24D0 CIRCLED LATIN SMALL LETTER A
	0x86C0: 'ⓑ' // U+24D1 CIRCLED LATIN SMALL LETTER B
	0x86C1: 'ⓒ' // U+24D2 CIRCLED LATIN SMALL LETTER C
	0x86C2: 'ⓓ' // U+24D3 CIRCLED LATIN SMALL LETTER D
	0x86C3: 'ⓔ' // U+24D4 CIRCLED LATIN SMALL LETTER E
	0x86C4: 'ⓕ' // U+24D5 CIRCLED LATIN SMALL LETTER F
	0x86C5: 'ⓖ' // U+24D6 CIRCLED LATIN SMALL LETTER G
	0x86C6: 'ⓗ' // U+24D7 CIRCLED LATIN SMALL LETTER H
	0x86C7: 'ⓘ' // U+24D8 CIRCLED LATIN SMALL LETTER I
	0x86C8: 'ⓙ' // U+24D9 CIRCLED LATIN SMALL LETTER J
	0x86C9: 'ⓚ' // U+24DA CIRCLED LATIN SMALL LETTER K
	0x86CA: 'ⓛ' // U+24DB CIRCLED LATIN SMALL LETTER L
	0x86CB: 'ⓜ' // U+24DC CIRCLED LATIN SMALL LETTER M
	0x86CC: 'ⓝ' // U+24DD CIRCLED LATIN SMALL LETTER N
	0x86CD: 'ⓞ' // U+24DE CIRCLED LATIN SMALL LETTER O
	0x86CE: 'ⓟ' // U+24DF CIRCLED LATIN SMALL LETTER P
	0x86CF: 'ⓠ' // U+24E0 CIRCLED LATIN SMALL LETTER Q
	0x86D0: 'ⓡ' // U+24E1 CIRCLED LATIN SMALL LETTER R
	0x86D1: 'ⓢ' // U+24E2 CIRCLED LATIN SMALL LETTER S
	0x86D2: 'ⓣ' // U+24E3 CIRCLED LATIN SMALL LETTER T
	0x86D3: 'ⓤ' // U+24E4 CIRCLED LATIN SMALL LETTER U
	0x86D4: 'ⓥ' // U+24E5 CIRCLED LATIN SMALL LETTER V
	0x86D5: 'ⓦ' // U+24E6 CIRCLED LATIN SMALL LETTER W
	0x86D6: 'ⓧ' // U+24E7 CIRCLED LATIN SMALL LETTER X
	0x86D7: 'ⓨ' // U+24E8 CIRCLED LATIN SMALL LETTER Y
	0x86D8: 'ⓩ' // U+24E9 CIRCLED LATIN SMALL LETTER Z
	0x86D9: '㋐' // U+32D0 CIRCLED KATAKANA A
	0x86DA: '㋑' // U+32D1 CIRCLED KATAKANA I
	0x86DB: '㋒' // U+32D2 CIRCLED KATAKANA U
	0x86DC: '㋓' // U+32D3 CIRCLED KATAKANA E
	0x86DD: '㋔' // U+32D4 CIRCLED KATAKANA O
	0x86DE: '㋕' // U+32D5 CIRCLED KATAKANA KA
	0x86DF: '㋖' // U+32D6 CIRCLED KATAKANA KI
	0x86E0: '㋗' // U+32D7 CIRCLED KATAKANA KU
	0x86E1: '㋘' // U+32D8 CIRCLED KATAKANA KE
	0x86E2: '㋙' // U+32D9 CIRCLED KATAKANA KO
	0x86E3: '㋚' // U+32DA CIRCLED KATAKANA SA
	0x86E4: '㋛' // U+32DB CIRCLED KATAKANA SI
	0x86E5: '㋜' // U+32DC CIRCLED KATAKANA SU
	0x86E6: '㋝' // U+32DD CIRCLED KATAKANA SE
	0x86E7: '㋞' // U+32DE CIRCLED KATAKANA SO
	0x86E8: '㋟' // U+32DF CIRCLED KATAKANA TA
	0x86E9: '㋠' // U+32E0 CIRCLED KATAKANA TI
	0x86EA: '㋡' // U+32E1 CIRCLED KATAKANA TU
	0x86EB: '㋢' // U+32E2 CIRCLED KATAKANA TE
	0x86EC: '㋣' // U+32E3 CIRCLED KATAKANA TO
	0x86ED: '㋺' // U+32FA CIRCLED KATAKANA RO
	0x86EE: '㋩' // U+32E9 CIRCLED KATAKANA HA
	0x86EF: '㋥' // U+32E5 CIRCLED KATAKANA NI
	0x86F0: '㋭' // U+32ED CIRCLED KATAKANA HO
	0x86F1: '㋬' // U+32EC CIRCLED KATAKANA HE
	0x86FB: '⁑' // U+2051 TWO ASTERISKS ALIGNED VERTICALLY
	0x86FC: '⁂' // U+2042 ASTERISM
	0x8740: '①' // U+2460 CIRCLED DIGIT ONE
	0x8741: '②' // U+2461 CIRCLED DIGIT TWO
	0x8742: '③' // U+2462 CIRCLED DIGIT THREE
	0x8743: '④' // U+2463 CIRCLED DIGIT FOUR
	0x8744: '⑤' // U+2464 CIRCLED DIGIT FIVE
	0x8745: '⑥' // U+2465 CIRCLED DIGIT SIX
	0x8746: '⑦' // U+2466 CIRCLED DIGIT SEVEN
	0x8747: '⑧' // U+2467 CIRCLED DIGIT EIGHT
	0x8748: '⑨' // U+2468 CIRCLED DIGIT NINE
	0x8749: '⑩' // U+2469 CIRCLED NUMBER TEN
	0x874A: '⑪' // U+246A CIRCLED NUMBER ELEVEN
	0x874B: '⑫' // U+246B CIRCLED NUMBER TWELVE
	0x874C: '⑬' // U+246C CIRCLED NUMBER THIRTEEN
	0x874D: '⑭' // U+246D CIRCLED NUMBER FOURTEEN
	0x874E: '⑮' // U+246E CIRCLED NUMBER FIFTEEN
	0x874F: '⑯' // U+246F CIRCLED NUMBER SIXTEEN
	0x8750: '⑰' // U+2470 CIRCLED NUMBER SEVENTEEN
	0x8751: '⑱' // U+2471 CIRCLED NUMBER EIGHTEEN
	0x8752: '⑲' // U+2472 CIRCLED NUMBER NINETEEN
	0x8753: '⑳' // U+2473 CIRCLED NUMBER TWENTY
	0x8754: 'Ⅰ' // U+2160 ROMAN NUMERAL ONE
	0x8755: 'Ⅱ' // U+2161 ROMAN NUMERAL TWO
	0x8756: 'Ⅲ' // U+2162 ROMAN NUMERAL THREE
	0x8757: 'Ⅳ' // U+2163 ROMAN NUMERAL FOUR
	0x8758: 'Ⅴ' // U+2164 ROMAN NUMERAL FIVE
	0x8759: 'Ⅵ' // U+2165 ROMAN NUMERAL SIX
	0x875A: 'Ⅶ' // U+2166 ROMAN NUMERAL SEVEN
	0x875B: 'Ⅷ' // U+2167 ROMAN NUMERAL EIGHT
	0x875C: 'Ⅸ' // U+2168 ROMAN NUMERAL NINE
	0x875D: 'Ⅹ' // U+2169 ROMAN NUMERAL TEN
	0x875E: 'Ⅺ' // U+216A ROMAN NUMERAL ELEVEN
	0x875F: '㍉' // U+3349 SQUARE MIRI
	0x8760: '㌔' // U+3314 SQUARE KIRO
	0x8761: '㌢' // U+3322 SQUARE SENTI
	0x8762: '㍍' // U+334D SQUARE MEETORU
	0x8763: '㌘' // U+3318 SQUARE GURAMU
	0x8764: '㌧' // U+3327 SQUARE TON
	0x8765: '㌃' // U+3303 SQUARE AARU
	0x8766: '㌶' // U+3336 SQUARE HEKUTAARU
	0x8767: '㍑' // U+3351 SQUARE RITTORU
	0x8768: '㍗' // U+3357 SQUARE WATTO
	0x8769: '㌍' // U+330D SQUARE KARORII
	0x876A: '㌦' // U+3326 SQUARE DORU
	0x876B: '㌣' // U+3323 SQUARE SENTO
	0x876C: '㌫' // U+332B SQUARE PAASENTO
	0x876D: '㍊' // U+334A SQUARE MIRIBAARU
	0x876E: '㌻' // U+333B SQUARE PEEZI
	0x876F: '㎜' // U+339C SQUARE MM
	0x8770: '㎝' // U+339D SQUARE CM
	0x8771: '㎞' // U+339E SQUARE KM
	0x8772: '㎎' // U+338E SQUARE MG
	0x8773: '㎏' // U+338F SQUARE KG
	0x8774: '㏄' // U+33C4 SQUARE CC
	0x8775: '㎡' // U+33A1 SQUARE M SQUARED
	0x8776: 'Ⅻ' // U+216B ROMAN NUMERAL TWELVE
	0x877E: '㍻' // U+337B SQUARE ERA NAME HEISEI
	0x8780: '〝' // U+301D REVERSED DOUBLE PRIME QUOTATION MARK
	0x8781: '〟' // U+301F LOW DOUBLE PRIME QUOTATION MARK
	0x8782: '№' // U+2116 NUMERO SIGN
	0x8783: '㏍' // U+33CD SQUARE KK
	0x8784: '℡' // U+2121 TELEPHONE SIGN
	0x8785: '㊤' // U+32A4 CIRCLED IDEOGRAPH HIGH
	0x8786: '㊥' // U+32A5 CIRCLED IDEOGRAPH CENTRE
	0x8787: '㊦' // U+32A6 CIRCLED IDEOGRAPH LOW
	0x8788: '㊧' // U+32A7 CIRCLED IDEOGRAPH LEFT
	0x8789: '㊨' // U+32A8 CIRCLED IDEOGRAPH RIGHT
	0x878A: '㈱' // U+3231 PARENTHESIZED IDEOGRAPH STOCK
	0x878B: '㈲' // U+3232 PARENTHESIZED IDEOGRAPH HAVE
	0x878C: '㈹' // U+3239 PARENTHESIZED IDEOGRAPH REPRESENT
	0x878D: '㍾' // U+337E SQUARE ERA NAME MEIZI
	0x878E: '㍽' // U+337D SQUARE ERA NAME TAISYOU
	0x878F: '㍼' // U+337C SQUARE ERA NAME SYOUWA
	0x8793: '∮' // U+222E CONTOUR INTEGRAL
	0x8798: '∟' // U+221F RIGHT ANGLE
	0x8799: '⊿' // U+22BF RIGHT TRIANGLE
	0x879D: '❖' // U+2756 BLACK DIAMOND MINUS WHITE X
	0x879E: '☞' // U+261E WHITE RIGHT POINTING INDEX
	0x879F: '俱' // U+4FF1 <cjk>
	0x87A0: '𠀋' // U+2000B <cjk>
	0x87A1: '㐂' // U+3402 <cjk>
	0x87A2: '丨' // U+4E28 <cjk>
	0x87A3: '丯' // U+4E2F <cjk>
	0x87A4: '丰' // U+4E30 <cjk>
	0x87A5: '亍' // U+4E8D <cjk>
	0x87A6: '仡' // U+4EE1 <cjk>
	0x87A7: '份' // U+4EFD <cjk>
	0x87A8: '仿' // U+4EFF <cjk>
	0x87A9: '伃' // U+4F03 <cjk>
	0x87AA: '伋' // U+4F0B <cjk>
	0x87AB: '你' // U+4F60 <cjk>
	0x87AC: '佈' // U+4F48 <cjk>
	0x87AD: '佉' // U+4F49 <cjk>
	0x87AE: '佖' // U+4F56 <cjk>
	0x87AF: '佟' // U+4F5F <cjk>
	0x87B0: '佪' // U+4F6A <cjk>
	0x87B1: '佬' // U+4F6C <cjk>
	0x87B2: '佾' // U+4F7E <cjk>
	0x87B3: '侊' // U+4F8A <cjk>
	0x87B4: '侔' // U+4F94 <cjk>
	0x87B5: '侗' // U+4F97 <cjk>
	0x87B6: '侮' // U+FA30 CJK COMPATIBILITY IDEOGRAPH-FA30
	0x87B7: '俉' // U+4FC9 <cjk>
	0x87B8: '俠' // U+4FE0 <cjk>
	0x87B9: '倁' // U+5001 <cjk>
	0x87BA: '倂' // U+5002 <cjk>
	0x87BB: '倎' // U+500E <cjk>
	0x87BC: '倘' // U+5018 <cjk>
	0x87BD: '倧' // U+5027 <cjk>
	0x87BE: '倮' // U+502E <cjk>
	0x87BF: '偀' // U+5040 <cjk>
	0x87C0: '倻' // U+503B <cjk>
	0x87C1: '偁' // U+5041 <cjk>
	0x87C2: '傔' // U+5094 <cjk>
	0x87C3: '僌' // U+50CC <cjk>
	0x87C4: '僲' // U+50F2 <cjk>
	0x87C5: '僐' // U+50D0 <cjk>
	0x87C6: '僦' // U+50E6 <cjk>
	0x87C7: '僧' // U+FA31 CJK COMPATIBILITY IDEOGRAPH-FA31
	0x87C8: '儆' // U+5106 <cjk>
	0x87C9: '儃' // U+5103 <cjk>
	0x87CA: '儋' // U+510B <cjk>
	0x87CB: '儞' // U+511E <cjk>
	0x87CC: '儵' // U+5135 <cjk>
	0x87CD: '兊' // U+514A <cjk>
	0x87CE: '免' // U+FA32 CJK COMPATIBILITY IDEOGRAPH-FA32
	0x87CF: '兕' // U+5155 <cjk>
	0x87D0: '兗' // U+5157 <cjk>
	0x87D1: '㒵' // U+34B5 <cjk>
	0x87D2: '冝' // U+519D <cjk>
	0x87D3: '凃' // U+51C3 <cjk>
	0x87D4: '凊' // U+51CA <cjk>
	0x87D5: '凞' // U+51DE <cjk>
	0x87D6: '凢' // U+51E2 <cjk>
	0x87D7: '凮' // U+51EE <cjk>
	0x87D8: '刁' // U+5201 <cjk>
	0x87D9: '㓛' // U+34DB <cjk>
	0x87DA: '刓' // U+5213 <cjk>
	0x87DB: '刕' // U+5215 <cjk>
	0x87DC: '剉' // U+5249 <cjk>
	0x87DD: '剗' // U+5257 <cjk>
	0x87DE: '剡' // U+5261 <cjk>
	0x87DF: '劓' // U+5293 <cjk>
	0x87E0: '勈' // U+52C8 <cjk>
	0x87E1: '勉' // U+FA33 CJK COMPATIBILITY IDEOGRAPH-FA33
	0x87E2: '勌' // U+52CC <cjk>
	0x87E3: '勐' // U+52D0 <cjk>
	0x87E4: '勖' // U+52D6 <cjk>
	0x87E5: '勛' // U+52DB <cjk>
	0x87E6: '勤' // U+FA34 CJK COMPATIBILITY IDEOGRAPH-FA34
	0x87E7: '勰' // U+52F0 <cjk>
	0x87E8: '勻' // U+52FB <cjk>
	0x87E9: '匀' // U+5300 <cjk>
	0x87EA: '匇' // U+5307 <cjk>
	0x87EB: '匜' // U+531C <cjk>
	0x87EC: '卑' // U+FA35 CJK COMPATIBILITY IDEOGRAPH-FA35
	0x87ED: '卡' // U+5361 <cjk>
	0x87EE: '卣' // U+5363 <cjk>
	0x87EF: '卽' // U+537D <cjk>
	0x87F0: '厓' // U+5393 <cjk>
	0x87F1: '厝' // U+539D <cjk>
	0x87F2: '厲' // U+53B2 <cjk>
	0x87F3: '吒' // U+5412 <cjk>
	0x87F4: '吧' // U+5427 <cjk>
	0x87F5: '呍' // U+544D <cjk>
	0x87F6: '咜' // U+549C <cjk>
	0x87F7: '呫' // U+546B <cjk>
	0x87F8: '呴' // U+5474 <cjk>
	0x87F9: '呿' // U+547F <cjk>
	0x87FA: '咈' // U+5488 <cjk>
	0x87FB: '咖' // U+5496 <cjk>
	0x87FC: '咡' // U+54A1 <cjk>
	0x8840: '咩' // U+54A9 <cjk>
	0x8841: '哆' // U+54C6 <cjk>
	0x8842: '哿' // U+54FF <cjk>
	0x8843: '唎' // U+550E <cjk>
	0x8844: '唫' // U+552B <cjk>
	0x8845: '唵' // U+5535 <cjk>
	0x8846: '啐' // U+5550 <cjk>
	0x8847: '啞' // U+555E <cjk>
	0x8848: '喁' // U+5581 <cjk>
	0x8849: '喆' // U+5586 <cjk>
	0x884A: '喎' // U+558E <cjk>
	0x884B: '喝' // U+FA36 CJK COMPATIBILITY IDEOGRAPH-FA36
	0x884C: '喭' // U+55AD <cjk>
	0x884D: '嗎' // U+55CE <cjk>
	0x884E: '嘆' // U+FA37 CJK COMPATIBILITY IDEOGRAPH-FA37
	0x884F: '嘈' // U+5608 <cjk>
	0x8850: '嘎' // U+560E <cjk>
	0x8851: '嘻' // U+563B <cjk>
	0x8852: '噉' // U+5649 <cjk>
	0x8853: '噶' // U+5676 <cjk>
	0x8854: '噦' // U+5666 <cjk>
	0x8855: '器' // U+FA38 CJK COMPATIBILITY IDEOGRAPH-FA38
	0x8856: '噯' // U+566F <cjk>
	0x8857: '噱' // U+5671 <cjk>
	0x8858: '噲' // U+5672 <cjk>
	0x8859: '嚙' // U+5699 <cjk>
	0x885A: '嚞' // U+569E <cjk>
	0x885B: '嚩' // U+56A9 <cjk>
	0x885C: '嚬' // U+56AC <cjk>
	0x885D: '嚳' // U+56B3 <cjk>
	0x885E: '囉' // U+56C9 <cjk>
	0x885F: '囊' // U+56CA <cjk>
	0x8860: '圊' // U+570A <cjk>
	0x8861: '𡈽' // U+2123D <cjk>
	0x8862: '圡' // U+5721 <cjk>
	0x8863: '圯' // U+572F <cjk>
	0x8864: '圳' // U+5733 <cjk>
	0x8865: '圴' // U+5734 <cjk>
	0x8866: '坰' // U+5770 <cjk>
	0x8867: '坷' // U+5777 <cjk>
	0x8868: '坼' // U+577C <cjk>
	0x8869: '垜' // U+579C <cjk>
	0x886A: '﨏' // U+FA0F CJK COMPATIBILITY IDEOGRAPH-FA0F
	0x886B: '𡌛' // U+2131B <cjk>
	0x886C: '垸' // U+57B8 <cjk>
	0x886D: '埇' // U+57C7 <cjk>
	0x886E: '埈' // U+57C8 <cjk>
	0x886F: '埏' // U+57CF <cjk>
	0x8870: '埤' // U+57E4 <cjk>
	0x8871: '埭' // U+57ED <cjk>
	0x8872: '埵' // U+57F5 <cjk>
	0x8873: '埶' // U+57F6 <cjk>
	0x8874: '埿' // U+57FF <cjk>
	0x8875: '堉' // U+5809 <cjk>
	0x8876: '塚' // U+FA10 CJK COMPATIBILITY IDEOGRAPH-FA10
	0x8877: '塡' // U+5861 <cjk>
	0x8878: '塤' // U+5864 <cjk>
	0x8879: '塀' // U+FA39 CJK COMPATIBILITY IDEOGRAPH-FA39
	0x887A: '塼' // U+587C <cjk>
	0x887B: '墉' // U+5889 <cjk>
	0x887C: '增' // U+589E <cjk>
	0x887D: '墨' // U+FA3A CJK COMPATIBILITY IDEOGRAPH-FA3A
	0x887E: '墩' // U+58A9 <cjk>
	0x8880: '𡑮' // U+2146E <cjk>
	0x8881: '壒' // U+58D2 <cjk>
	0x8882: '壎' // U+58CE <cjk>
	0x8883: '壔' // U+58D4 <cjk>
	0x8884: '壚' // U+58DA <cjk>
	0x8885: '壠' // U+58E0 <cjk>
	0x8886: '壩' // U+58E9 <cjk>
	0x8887: '夌' // U+590C <cjk>
	0x8888: '虁' // U+8641 <cjk>
	0x8889: '奝' // U+595D <cjk>
	0x888A: '奭' // U+596D <cjk>
	0x888B: '妋' // U+598B <cjk>
	0x888C: '妒' // U+5992 <cjk>
	0x888D: '妤' // U+59A4 <cjk>
	0x888E: '姃' // U+59C3 <cjk>
	0x888F: '姒' // U+59D2 <cjk>
	0x8890: '姝' // U+59DD <cjk>
	0x8891: '娓' // U+5A13 <cjk>
	0x8892: '娣' // U+5A23 <cjk>
	0x8893: '婧' // U+5A67 <cjk>
	0x8894: '婭' // U+5A6D <cjk>
	0x8895: '婷' // U+5A77 <cjk>
	0x8896: '婾' // U+5A7E <cjk>
	0x8897: '媄' // U+5A84 <cjk>
	0x8898: '媞' // U+5A9E <cjk>
	0x8899: '媧' // U+5AA7 <cjk>
	0x889A: '嫄' // U+5AC4 <cjk>
	0x889B: '𡢽' // U+218BD <cjk>
	0x889C: '嬙' // U+5B19 <cjk>
	0x889D: '嬥' // U+5B25 <cjk>
	0x889E: '剝' // U+525D <cjk>
	0x889F: '亜' // U+4E9C <cjk>
	0x88A0: '唖' // U+5516 <cjk>
	0x88A1: '娃' // U+5A03 <cjk>
	0x88A2: '阿' // U+963F <cjk>
	0x88A3: '哀' // U+54C0 <cjk>
	0x88A4: '愛' // U+611B <cjk>
	0x88A5: '挨' // U+6328 <cjk>
	0x88A6: '姶' // U+59F6 <cjk>
	0x88A7: '逢' // U+9022 <cjk>
	0x88A8: '葵' // U+8475 <cjk>
	0x88A9: '茜' // U+831C <cjk>
	0x88AA: '穐' // U+7A50 <cjk>
	0x88AB: '悪' // U+60AA <cjk>
	0x88AC: '握' // U+63E1 <cjk>
	0x88AD: '渥' // U+6E25 <cjk>
	0x88AE: '旭' // U+65ED <cjk>
	0x88AF: '葦' // U+8466 <cjk>
	0x88B0: '芦' // U+82A6 <cjk>
	0x88B1: '鯵' // U+9BF5 <cjk>
	0x88B2: '梓' // U+6893 <cjk>
	0x88B3: '圧' // U+5727 <cjk>
	0x88B4: '斡' // U+65A1 <cjk>
	0x88B5: '扱' // U+6271 <cjk>
	0x88B6: '宛' // U+5B9B <cjk>
	0x88B7: '姐' // U+59D0 <cjk>
	0x88B8: '虻' // U+867B <cjk>
	0x88B9: '飴' // U+98F4 <cjk>
	0x88BA: '絢' // U+7D62 <cjk>
	0x88BB: '綾' // U+7DBE <cjk>
	0x88BC: '鮎' // U+9B8E <cjk>
	0x88BD: '或' // U+6216 <cjk>
	0x88BE: '粟' // U+7C9F <cjk>
	0x88BF: '袷' // U+88B7 <cjk>
	0x88C0: '安' // U+5B89 <cjk>
	0x88C1: '庵' // U+5EB5 <cjk>
	0x88C2: '按' // U+6309 <cjk>
	0x88C3: '暗' // U+6697 <cjk>
	0x88C4: '案' // U+6848 <cjk>
	0x88C5: '闇' // U+95C7 <cjk>
	0x88C6: '鞍' // U+978D <cjk>
	0x88C7: '杏' // U+674F <cjk>
	0x88C8: '以' // U+4EE5 <cjk>
	0x88C9: '伊' // U+4F0A <cjk>
	0x88CA: '位' // U+4F4D <cjk>
	0x88CB: '依' // U+4F9D <cjk>
	0x88CC: '偉' // U+5049 <cjk>
	0x88CD: '囲' // U+56F2 <cjk>
	0x88CE: '夷' // U+5937 <cjk>
	0x88CF: '委' // U+59D4 <cjk>
	0x88D0: '威' // U+5A01 <cjk>
	0x88D1: '尉' // U+5C09 <cjk>
	0x88D2: '惟' // U+60DF <cjk>
	0x88D3: '意' // U+610F <cjk>
	0x88D4: '慰' // U+6170 <cjk>
	0x88D5: '易' // U+6613 <cjk>
	0x88D6: '椅' // U+6905 <cjk>
	0x88D7: '為' // U+70BA <cjk>
	0x88D8: '畏' // U+754F <cjk>
	0x88D9: '異' // U+7570 <cjk>
	0x88DA: '移' // U+79FB <cjk>
	0x88DB: '維' // U+7DAD <cjk>
	0x88DC: '緯' // U+7DEF <cjk>
	0x88DD: '胃' // U+80C3 <cjk>
	0x88DE: '萎' // U+840E <cjk>
	0x88DF: '衣' // U+8863 <cjk>
	0x88E0: '謂' // U+8B02 <cjk>
	0x88E1: '違' // U+9055 <cjk>
	0x88E2: '遺' // U+907A <cjk>
	0x88E3: '医' // U+533B <cjk>
	0x88E4: '井' // U+4E95 <cjk>
	0x88E5: '亥' // U+4EA5 <cjk>
	0x88E6: '域' // U+57DF <cjk>
	0x88E7: '育' // U+80B2 <cjk>
	0x88E8: '郁' // U+90C1 <cjk>
	0x88E9: '磯' // U+78EF <cjk>
	0x88EA: '一' // U+4E00 <cjk>
	0x88EB: '壱' // U+58F1 <cjk>
	0x88EC: '溢' // U+6EA2 <cjk>
	0x88ED: '逸' // U+9038 <cjk>
	0x88EE: '稲' // U+7A32 <cjk>
	0x88EF: '茨' // U+8328 <cjk>
	0x88F0: '芋' // U+828B <cjk>
	0x88F1: '鰯' // U+9C2F <cjk>
	0x88F2: '允' // U+5141 <cjk>
	0x88F3: '印' // U+5370 <cjk>
	0x88F4: '咽' // U+54BD <cjk>
	0x88F5: '員' // U+54E1 <cjk>
	0x88F6: '因' // U+56E0 <cjk>
	0x88F7: '姻' // U+59FB <cjk>
	0x88F8: '引' // U+5F15 <cjk>
	0x88F9: '飲' // U+98F2 <cjk>
	0x88FA: '淫' // U+6DEB <cjk>
	0x88FB: '胤' // U+80E4 <cjk>
	0x88FC: '蔭' // U+852D <cjk>
	0x8940: '院' // U+9662 <cjk>
	0x8941: '陰' // U+9670 <cjk>
	0x8942: '隠' // U+96A0 <cjk>
	0x8943: '韻' // U+97FB <cjk>
	0x8944: '吋' // U+540B <cjk>
	0x8945: '右' // U+53F3 <cjk>
	0x8946: '宇' // U+5B87 <cjk>
	0x8947: '烏' // U+70CF <cjk>
	0x8948: '羽' // U+7FBD <cjk>
	0x8949: '迂' // U+8FC2 <cjk>
	0x894A: '雨' // U+96E8 <cjk>
	0x894B: '卯' // U+536F <cjk>
	0x894C: '鵜' // U+9D5C <cjk>
	0x894D: '窺' // U+7ABA <cjk>
	0x894E: '丑' // U+4E11 <cjk>
	0x894F: '碓' // U+7893 <cjk>
	0x8950: '臼' // U+81FC <cjk>
	0x8951: '渦' // U+6E26 <cjk>
	0x8952: '嘘' // U+5618 <cjk>
	0x8953: '唄' // U+5504 <cjk>
	0x8954: '欝' // U+6B1D <cjk>
	0x8955: '蔚' // U+851A <cjk>
	0x8956: '鰻' // U+9C3B <cjk>
	0x8957: '姥' // U+59E5 <cjk>
	0x8958: '厩' // U+53A9 <cjk>
	0x8959: '浦' // U+6D66 <cjk>
	0x895A: '瓜' // U+74DC <cjk>
	0x895B: '閏' // U+958F <cjk>
	0x895C: '噂' // U+5642 <cjk>
	0x895D: '云' // U+4E91 <cjk>
	0x895E: '運' // U+904B <cjk>
	0x895F: '雲' // U+96F2 <cjk>
	0x8960: '荏' // U+834F <cjk>
	0x8961: '餌' // U+990C <cjk>
	0x8962: '叡' // U+53E1 <cjk>
	0x8963: '営' // U+55B6 <cjk>
	0x8964: '嬰' // U+5B30 <cjk>
	0x8965: '影' // U+5F71 <cjk>
	0x8966: '映' // U+6620 <cjk>
	0x8967: '曳' // U+66F3 <cjk>
	0x8968: '栄' // U+6804 <cjk>
	0x8969: '永' // U+6C38 <cjk>
	0x896A: '泳' // U+6CF3 <cjk>
	0x896B: '洩' // U+6D29 <cjk>
	0x896C: '瑛' // U+745B <cjk>
	0x896D: '盈' // U+76C8 <cjk>
	0x896E: '穎' // U+7A4E <cjk>
	0x896F: '頴' // U+9834 <cjk>
	0x8970: '英' // U+82F1 <cjk>
	0x8971: '衛' // U+885B <cjk>
	0x8972: '詠' // U+8A60 <cjk>
	0x8973: '鋭' // U+92ED <cjk>
	0x8974: '液' // U+6DB2 <cjk>
	0x8975: '疫' // U+75AB <cjk>
	0x8976: '益' // U+76CA <cjk>
	0x8977: '駅' // U+99C5 <cjk>
	0x8978: '悦' // U+60A6 <cjk>
	0x8979: '謁' // U+8B01 <cjk>
	0x897A: '越' // U+8D8A <cjk>
	0x897B: '閲' // U+95B2 <cjk>
	0x897C: '榎' // U+698E <cjk>
	0x897D: '厭' // U+53AD <cjk>
	0x897E: '円' // U+5186 <cjk>
	0x8980: '園' // U+5712 <cjk>
	0x8981: '堰' // U+5830 <cjk>
	0x8982: '奄' // U+5944 <cjk>
	0x8983: '宴' // U+5BB4 <cjk>
	0x8984: '延' // U+5EF6 <cjk>
	0x8985: '怨' // U+6028 <cjk>
	0x8986: '掩' // U+63A9 <cjk>
	0x8987: '援' // U+63F4 <cjk>
	0x8988: '沿' // U+6CBF <cjk>
	0x8989: '演' // U+6F14 <cjk>
	0x898A: '炎' // U+708E <cjk>
	0x898B: '焔' // U+7114 <cjk>
	0x898C: '煙' // U+7159 <cjk>
	0x898D: '燕' // U+71D5 <cjk>
	0x898E: '猿' // U+733F <cjk>
	0x898F: '縁' // U+7E01 <cjk>
	0x8990: '艶' // U+8276 <cjk>
	0x8991: '苑' // U+82D1 <cjk>
	0x8992: '薗' // U+8597 <cjk>
	0x8993: '遠' // U+9060 <cjk>
	0x8994: '鉛' // U+925B <cjk>
	0x8995: '鴛' // U+9D1B <cjk>
	0x8996: '塩' // U+5869 <cjk>
	0x8997: '於' // U+65BC <cjk>
	0x8998: '汚' // U+6C5A <cjk>
	0x8999: '甥' // U+7525 <cjk>
	0x899A: '凹' // U+51F9 <cjk>
	0x899B: '央' // U+592E <cjk>
	0x899C: '奥' // U+5965 <cjk>
	0x899D: '往' // U+5F80 <cjk>
	0x899E: '応' // U+5FDC <cjk>
	0x899F: '押' // U+62BC <cjk>
	0x89A0: '旺' // U+65FA <cjk>
	0x89A1: '横' // U+6A2A <cjk>
	0x89A2: '欧' // U+6B27 <cjk>
	0x89A3: '殴' // U+6BB4 <cjk>
	0x89A4: '王' // U+738B <cjk>
	0x89A5: '翁' // U+7FC1 <cjk>
	0x89A6: '襖' // U+8956 <cjk>
	0x89A7: '鴬' // U+9D2C <cjk>
	0x89A8: '鴎' // U+9D0E <cjk>
	0x89A9: '黄' // U+9EC4 <cjk>
	0x89AA: '岡' // U+5CA1 <cjk>
	0x89AB: '沖' // U+6C96 <cjk>
	0x89AC: '荻' // U+837B <cjk>
	0x89AD: '億' // U+5104 <cjk>
	0x89AE: '屋' // U+5C4B <cjk>
	0x89AF: '憶' // U+61B6 <cjk>
	0x89B0: '臆' // U+81C6 <cjk>
	0x89B1: '桶' // U+6876 <cjk>
	0x89B2: '牡' // U+7261 <cjk>
	0x89B3: '乙' // U+4E59 <cjk>
	0x89B4: '俺' // U+4FFA <cjk>
	0x89B5: '卸' // U+5378 <cjk>
	0x89B6: '恩' // U+6069 <cjk>
	0x89B7: '温' // U+6E29 <cjk>
	0x89B8: '穏' // U+7A4F <cjk>
	0x89B9: '音' // U+97F3 <cjk>
	0x89BA: '下' // U+4E0B <cjk>
	0x89BB: '化' // U+5316 <cjk>
	0x89BC: '仮' // U+4EEE <cjk>
	0x89BD: '何' // U+4F55 <cjk>
	0x89BE: '伽' // U+4F3D <cjk>
	0x89BF: '価' // U+4FA1 <cjk>
	0x89C0: '佳' // U+4F73 <cjk>
	0x89C1: '加' // U+52A0 <cjk>
	0x89C2: '可' // U+53EF <cjk>
	0x89C3: '嘉' // U+5609 <cjk>
	0x89C4: '夏' // U+590F <cjk>
	0x89C5: '嫁' // U+5AC1 <cjk>
	0x89C6: '家' // U+5BB6 <cjk>
	0x89C7: '寡' // U+5BE1 <cjk>
	0x89C8: '科' // U+79D1 <cjk>
	0x89C9: '暇' // U+6687 <cjk>
	0x89CA: '果' // U+679C <cjk>
	0x89CB: '架' // U+67B6 <cjk>
	0x89CC: '歌' // U+6B4C <cjk>
	0x89CD: '河' // U+6CB3 <cjk>
	0x89CE: '火' // U+706B <cjk>
	0x89CF: '珂' // U+73C2 <cjk>
	0x89D0: '禍' // U+798D <cjk>
	0x89D1: '禾' // U+79BE <cjk>
	0x89D2: '稼' // U+7A3C <cjk>
	0x89D3: '箇' // U+7B87 <cjk>
	0x89D4: '花' // U+82B1 <cjk>
	0x89D5: '苛' // U+82DB <cjk>
	0x89D6: '茄' // U+8304 <cjk>
	0x89D7: '荷' // U+8377 <cjk>
	0x89D8: '華' // U+83EF <cjk>
	0x89D9: '菓' // U+83D3 <cjk>
	0x89DA: '蝦' // U+8766 <cjk>
	0x89DB: '課' // U+8AB2 <cjk>
	0x89DC: '嘩' // U+5629 <cjk>
	0x89DD: '貨' // U+8CA8 <cjk>
	0x89DE: '迦' // U+8FE6 <cjk>
	0x89DF: '過' // U+904E <cjk>
	0x89E0: '霞' // U+971E <cjk>
	0x89E1: '蚊' // U+868A <cjk>
	0x89E2: '俄' // U+4FC4 <cjk>
	0x89E3: '峨' // U+5CE8 <cjk>
	0x89E4: '我' // U+6211 <cjk>
	0x89E5: '牙' // U+7259 <cjk>
	0x89E6: '画' // U+753B <cjk>
	0x89E7: '臥' // U+81E5 <cjk>
	0x89E8: '芽' // U+82BD <cjk>
	0x89E9: '蛾' // U+86FE <cjk>
	0x89EA: '賀' // U+8CC0 <cjk>
	0x89EB: '雅' // U+96C5 <cjk>
	0x89EC: '餓' // U+9913 <cjk>
	0x89ED: '駕' // U+99D5 <cjk>
	0x89EE: '介' // U+4ECB <cjk>
	0x89EF: '会' // U+4F1A <cjk>
	0x89F0: '解' // U+89E3 <cjk>
	0x89F1: '回' // U+56DE <cjk>
	0x89F2: '塊' // U+584A <cjk>
	0x89F3: '壊' // U+58CA <cjk>
	0x89F4: '廻' // U+5EFB <cjk>
	0x89F5: '快' // U+5FEB <cjk>
	0x89F6: '怪' // U+602A <cjk>
	0x89F7: '悔' // U+6094 <cjk>
	0x89F8: '恢' // U+6062 <cjk>
	0x89F9: '懐' // U+61D0 <cjk>
	0x89FA: '戒' // U+6212 <cjk>
	0x89FB: '拐' // U+62D0 <cjk>
	0x89FC: '改' // U+6539 <cjk>
	0x8A40: '魁' // U+9B41 <cjk>
	0x8A41: '晦' // U+6666 <cjk>
	0x8A42: '械' // U+68B0 <cjk>
	0x8A43: '海' // U+6D77 <cjk>
	0x8A44: '灰' // U+7070 <cjk>
	0x8A45: '界' // U+754C <cjk>
	0x8A46: '皆' // U+7686 <cjk>
	0x8A47: '絵' // U+7D75 <cjk>
	0x8A48: '芥' // U+82A5 <cjk>
	0x8A49: '蟹' // U+87F9 <cjk>
	0x8A4A: '開' // U+958B <cjk>
	0x8A4B: '階' // U+968E <cjk>
	0x8A4C: '貝' // U+8C9D <cjk>
	0x8A4D: '凱' // U+51F1 <cjk>
	0x8A4E: '劾' // U+52BE <cjk>
	0x8A4F: '外' // U+5916 <cjk>
	0x8A50: '咳' // U+54B3 <cjk>
	0x8A51: '害' // U+5BB3 <cjk>
	0x8A52: '崖' // U+5D16 <cjk>
	0x8A53: '慨' // U+6168 <cjk>
	0x8A54: '概' // U+6982 <cjk>
	0x8A55: '涯' // U+6DAF <cjk>
	0x8A56: '碍' // U+788D <cjk>
	0x8A57: '蓋' // U+84CB <cjk>
	0x8A58: '街' // U+8857 <cjk>
	0x8A59: '該' // U+8A72 <cjk>
	0x8A5A: '鎧' // U+93A7 <cjk>
	0x8A5B: '骸' // U+9AB8 <cjk>
	0x8A5C: '浬' // U+6D6C <cjk>
	0x8A5D: '馨' // U+99A8 <cjk>
	0x8A5E: '蛙' // U+86D9 <cjk>
	0x8A5F: '垣' // U+57A3 <cjk>
	0x8A60: '柿' // U+67FF <cjk>
	0x8A61: '蛎' // U+86CE <cjk>
	0x8A62: '鈎' // U+920E <cjk>
	0x8A63: '劃' // U+5283 <cjk>
	0x8A64: '嚇' // U+5687 <cjk>
	0x8A65: '各' // U+5404 <cjk>
	0x8A66: '廓' // U+5ED3 <cjk>
	0x8A67: '拡' // U+62E1 <cjk>
	0x8A68: '撹' // U+64B9 <cjk>
	0x8A69: '格' // U+683C <cjk>
	0x8A6A: '核' // U+6838 <cjk>
	0x8A6B: '殻' // U+6BBB <cjk>
	0x8A6C: '獲' // U+7372 <cjk>
	0x8A6D: '確' // U+78BA <cjk>
	0x8A6E: '穫' // U+7A6B <cjk>
	0x8A6F: '覚' // U+899A <cjk>
	0x8A70: '角' // U+89D2 <cjk>
	0x8A71: '赫' // U+8D6B <cjk>
	0x8A72: '較' // U+8F03 <cjk>
	0x8A73: '郭' // U+90ED <cjk>
	0x8A74: '閣' // U+95A3 <cjk>
	0x8A75: '隔' // U+9694 <cjk>
	0x8A76: '革' // U+9769 <cjk>
	0x8A77: '学' // U+5B66 <cjk>
	0x8A78: '岳' // U+5CB3 <cjk>
	0x8A79: '楽' // U+697D <cjk>
	0x8A7A: '額' // U+984D <cjk>
	0x8A7B: '顎' // U+984E <cjk>
	0x8A7C: '掛' // U+639B <cjk>
	0x8A7D: '笠' // U+7B20 <cjk>
	0x8A7E: '樫' // U+6A2B <cjk>
	0x8A80: '橿' // U+6A7F <cjk>
	0x8A81: '梶' // U+68B6 <cjk>
	0x8A82: '鰍' // U+9C0D <cjk>
	0x8A83: '潟' // U+6F5F <cjk>
	0x8A84: '割' // U+5272 <cjk>
	0x8A85: '喝' // U+559D <cjk>
	0x8A86: '恰' // U+6070 <cjk>
	0x8A87: '括' // U+62EC <cjk>
	0x8A88: '活' // U+6D3B <cjk>
	0x8A89: '渇' // U+6E07 <cjk>
	0x8A8A: '滑' // U+6ED1 <cjk>
	0x8A8B: '葛' // U+845B <cjk>
	0x8A8C: '褐' // U+8910 <cjk>
	0x8A8D: '轄' // U+8F44 <cjk>
	0x8A8E: '且' // U+4E14 <cjk>
	0x8A8F: '鰹' // U+9C39 <cjk>
	0x8A90: '叶' // U+53F6 <cjk>
	0x8A91: '椛' // U+691B <cjk>
	0x8A92: '樺' // U+6A3A <cjk>
	0x8A93: '鞄' // U+9784 <cjk>
	0x8A94: '株' // U+682A <cjk>
	0x8A95: '兜' // U+515C <cjk>
	0x8A96: '竃' // U+7AC3 <cjk>
	0x8A97: '蒲' // U+84B2 <cjk>
	0x8A98: '釜' // U+91DC <cjk>
	0x8A99: '鎌' // U+938C <cjk>
	0x8A9A: '噛' // U+565B <cjk>
	0x8A9B: '鴨' // U+9D28 <cjk>
	0x8A9C: '栢' // U+6822 <cjk>
	0x8A9D: '茅' // U+8305 <cjk>
	0x8A9E: '萱' // U+8431 <cjk>
	0x8A9F: '粥' // U+7CA5 <cjk>
	0x8AA0: '刈' // U+5208 <cjk>
	0x8AA1: '苅' // U+82C5 <cjk>
	0x8AA2: '瓦' // U+74E6 <cjk>
	0x8AA3: '乾' // U+4E7E <cjk>
	0x8AA4: '侃' // U+4F83 <cjk>
	0x8AA5: '冠' // U+51A0 <cjk>
	0x8AA6: '寒' // U+5BD2 <cjk>
	0x8AA7: '刊' // U+520A <cjk>
	0x8AA8: '勘' // U+52D8 <cjk>
	0x8AA9: '勧' // U+52E7 <cjk>
	0x8AAA: '巻' // U+5DFB <cjk>
	0x8AAB: '喚' // U+559A <cjk>
	0x8AAC: '堪' // U+582A <cjk>
	0x8AAD: '姦' // U+59E6 <cjk>
	0x8AAE: '完' // U+5B8C <cjk>
	0x8AAF: '官' // U+5B98 <cjk>
	0x8AB0: '寛' // U+5BDB <cjk>
	0x8AB1: '干' // U+5E72 <cjk>
	0x8AB2: '幹' // U+5E79 <cjk>
	0x8AB3: '患' // U+60A3 <cjk>
	0x8AB4: '感' // U+611F <cjk>
	0x8AB5: '慣' // U+6163 <cjk>
	0x8AB6: '憾' // U+61BE <cjk>
	0x8AB7: '換' // U+63DB <cjk>
	0x8AB8: '敢' // U+6562 <cjk>
	0x8AB9: '柑' // U+67D1 <cjk>
	0x8ABA: '桓' // U+6853 <cjk>
	0x8ABB: '棺' // U+68FA <cjk>
	0x8ABC: '款' // U+6B3E <cjk>
	0x8ABD: '歓' // U+6B53 <cjk>
	0x8ABE: '汗' // U+6C57 <cjk>
	0x8ABF: '漢' // U+6F22 <cjk>
	0x8AC0: '澗' // U+6F97 <cjk>
	0x8AC1: '潅' // U+6F45 <cjk>
	0x8AC2: '環' // U+74B0 <cjk>
	0x8AC3: '甘' // U+7518 <cjk>
	0x8AC4: '監' // U+76E3 <cjk>
	0x8AC5: '看' // U+770B <cjk>
	0x8AC6: '竿' // U+7AFF <cjk>
	0x8AC7: '管' // U+7BA1 <cjk>
	0x8AC8: '簡' // U+7C21 <cjk>
	0x8AC9: '緩' // U+7DE9 <cjk>
	0x8ACA: '缶' // U+7F36 <cjk>
	0x8ACB: '翰' // U+7FF0 <cjk>
	0x8ACC: '肝' // U+809D <cjk>
	0x8ACD: '艦' // U+8266 <cjk>
	0x8ACE: '莞' // U+839E <cjk>
	0x8ACF: '観' // U+89B3 <cjk>
	0x8AD0: '諌' // U+8ACC <cjk>
	0x8AD1: '貫' // U+8CAB <cjk>
	0x8AD2: '還' // U+9084 <cjk>
	0x8AD3: '鑑' // U+9451 <cjk>
	0x8AD4: '間' // U+9593 <cjk>
	0x8AD5: '閑' // U+9591 <cjk>
	0x8AD6: '関' // U+95A2 <cjk>
	0x8AD7: '陥' // U+9665 <cjk>
	0x8AD8: '韓' // U+97D3 <cjk>
	0x8AD9: '館' // U+9928 <cjk>
	0x8ADA: '舘' // U+8218 <cjk>
	0x8ADB: '丸' // U+4E38 <cjk>
	0x8ADC: '含' // U+542B <cjk>
	0x8ADD: '岸' // U+5CB8 <cjk>
	0x8ADE: '巌' // U+5DCC <cjk>
	0x8ADF: '玩' // U+73A9 <cjk>
	0x8AE0: '癌' // U+764C <cjk>
	0x8AE1: '眼' // U+773C <cjk>
	0x8AE2: '岩' // U+5CA9 <cjk>
	0x8AE3: '翫' // U+7FEB <cjk>
	0x8AE4: '贋' // U+8D0B <cjk>
	0x8AE5: '雁' // U+96C1 <cjk>
	0x8AE6: '頑' // U+9811 <cjk>
	0x8AE7: '顔' // U+9854 <cjk>
	0x8AE8: '願' // U+9858 <cjk>
	0x8AE9: '企' // U+4F01 <cjk>
	0x8AEA: '伎' // U+4F0E <cjk>
	0x8AEB: '危' // U+5371 <cjk>
	0x8AEC: '喜' // U+559C <cjk>
	0x8AED: '器' // U+5668 <cjk>
	0x8AEE: '基' // U+57FA <cjk>
	0x8AEF: '奇' // U+5947 <cjk>
	0x8AF0: '嬉' // U+5B09 <cjk>
	0x8AF1: '寄' // U+5BC4 <cjk>
	0x8AF2: '岐' // U+5C90 <cjk>
	0x8AF3: '希' // U+5E0C <cjk>
	0x8AF4: '幾' // U+5E7E <cjk>
	0x8AF5: '忌' // U+5FCC <cjk>
	0x8AF6: '揮' // U+63EE <cjk>
	0x8AF7: '机' // U+673A <cjk>
	0x8AF8: '旗' // U+65D7 <cjk>
	0x8AF9: '既' // U+65E2 <cjk>
	0x8AFA: '期' // U+671F <cjk>
	0x8AFB: '棋' // U+68CB <cjk>
	0x8AFC: '棄' // U+68C4 <cjk>
	0x8B40: '機' // U+6A5F <cjk>
	0x8B41: '帰' // U+5E30 <cjk>
	0x8B42: '毅' // U+6BC5 <cjk>
	0x8B43: '気' // U+6C17 <cjk>
	0x8B44: '汽' // U+6C7D <cjk>
	0x8B45: '畿' // U+757F <cjk>
	0x8B46: '祈' // U+7948 <cjk>
	0x8B47: '季' // U+5B63 <cjk>
	0x8B48: '稀' // U+7A00 <cjk>
	0x8B49: '紀' // U+7D00 <cjk>
	0x8B4A: '徽' // U+5FBD <cjk>
	0x8B4B: '規' // U+898F <cjk>
	0x8B4C: '記' // U+8A18 <cjk>
	0x8B4D: '貴' // U+8CB4 <cjk>
	0x8B4E: '起' // U+8D77 <cjk>
	0x8B4F: '軌' // U+8ECC <cjk>
	0x8B50: '輝' // U+8F1D <cjk>
	0x8B51: '飢' // U+98E2 <cjk>
	0x8B52: '騎' // U+9A0E <cjk>
	0x8B53: '鬼' // U+9B3C <cjk>
	0x8B54: '亀' // U+4E80 <cjk>
	0x8B55: '偽' // U+507D <cjk>
	0x8B56: '儀' // U+5100 <cjk>
	0x8B57: '妓' // U+5993 <cjk>
	0x8B58: '宜' // U+5B9C <cjk>
	0x8B59: '戯' // U+622F <cjk>
	0x8B5A: '技' // U+6280 <cjk>
	0x8B5B: '擬' // U+64EC <cjk>
	0x8B5C: '欺' // U+6B3A <cjk>
	0x8B5D: '犠' // U+72A0 <cjk>
	0x8B5E: '疑' // U+7591 <cjk>
	0x8B5F: '祇' // U+7947 <cjk>
	0x8B60: '義' // U+7FA9 <cjk>
	0x8B61: '蟻' // U+87FB <cjk>
	0x8B62: '誼' // U+8ABC <cjk>
	0x8B63: '議' // U+8B70 <cjk>
	0x8B64: '掬' // U+63AC <cjk>
	0x8B65: '菊' // U+83CA <cjk>
	0x8B66: '鞠' // U+97A0 <cjk>
	0x8B67: '吉' // U+5409 <cjk>
	0x8B68: '吃' // U+5403 <cjk>
	0x8B69: '喫' // U+55AB <cjk>
	0x8B6A: '桔' // U+6854 <cjk>
	0x8B6B: '橘' // U+6A58 <cjk>
	0x8B6C: '詰' // U+8A70 <cjk>
	0x8B6D: '砧' // U+7827 <cjk>
	0x8B6E: '杵' // U+6775 <cjk>
	0x8B6F: '黍' // U+9ECD <cjk>
	0x8B70: '却' // U+5374 <cjk>
	0x8B71: '客' // U+5BA2 <cjk>
	0x8B72: '脚' // U+811A <cjk>
	0x8B73: '虐' // U+8650 <cjk>
	0x8B74: '逆' // U+9006 <cjk>
	0x8B75: '丘' // U+4E18 <cjk>
	0x8B76: '久' // U+4E45 <cjk>
	0x8B77: '仇' // U+4EC7 <cjk>
	0x8B78: '休' // U+4F11 <cjk>
	0x8B79: '及' // U+53CA <cjk>
	0x8B7A: '吸' // U+5438 <cjk>
	0x8B7B: '宮' // U+5BAE <cjk>
	0x8B7C: '弓' // U+5F13 <cjk>
	0x8B7D: '急' // U+6025 <cjk>
	0x8B7E: '救' // U+6551 <cjk>
	0x8B80: '朽' // U+673D <cjk>
	0x8B81: '求' // U+6C42 <cjk>
	0x8B82: '汲' // U+6C72 <cjk>
	0x8B83: '泣' // U+6CE3 <cjk>
	0x8B84: '灸' // U+7078 <cjk>
	0x8B85: '球' // U+7403 <cjk>
	0x8B86: '究' // U+7A76 <cjk>
	0x8B87: '窮' // U+7AAE <cjk>
	0x8B88: '笈' // U+7B08 <cjk>
	0x8B89: '級' // U+7D1A <cjk>
	0x8B8A: '糾' // U+7CFE <cjk>
	0x8B8B: '給' // U+7D66 <cjk>
	0x8B8C: '旧' // U+65E7 <cjk>
	0x8B8D: '牛' // U+725B <cjk>
	0x8B8E: '去' // U+53BB <cjk>
	0x8B8F: '居' // U+5C45 <cjk>
	0x8B90: '巨' // U+5DE8 <cjk>
	0x8B91: '拒' // U+62D2 <cjk>
	0x8B92: '拠' // U+62E0 <cjk>
	0x8B93: '挙' // U+6319 <cjk>
	0x8B94: '渠' // U+6E20 <cjk>
	0x8B95: '虚' // U+865A <cjk>
	0x8B96: '許' // U+8A31 <cjk>
	0x8B97: '距' // U+8DDD <cjk>
	0x8B98: '鋸' // U+92F8 <cjk>
	0x8B99: '漁' // U+6F01 <cjk>
	0x8B9A: '禦' // U+79A6 <cjk>
	0x8B9B: '魚' // U+9B5A <cjk>
	0x8B9C: '亨' // U+4EA8 <cjk>
	0x8B9D: '享' // U+4EAB <cjk>
	0x8B9E: '京' // U+4EAC <cjk>
	0x8B9F: '供' // U+4F9B <cjk>
	0x8BA0: '侠' // U+4FA0 <cjk>
	0x8BA1: '僑' // U+50D1 <cjk>
	0x8BA2: '兇' // U+5147 <cjk>
	0x8BA3: '競' // U+7AF6 <cjk>
	0x8BA4: '共' // U+5171 <cjk>
	0x8BA5: '凶' // U+51F6 <cjk>
	0x8BA6: '協' // U+5354 <cjk>
	0x8BA7: '匡' // U+5321 <cjk>
	0x8BA8: '卿' // U+537F <cjk>
	0x8BA9: '叫' // U+53EB <cjk>
	0x8BAA: '喬' // U+55AC <cjk>
	0x8BAB: '境' // U+5883 <cjk>
	0x8BAC: '峡' // U+5CE1 <cjk>
	0x8BAD: '強' // U+5F37 <cjk>
	0x8BAE: '彊' // U+5F4A <cjk>
	0x8BAF: '怯' // U+602F <cjk>
	0x8BB0: '恐' // U+6050 <cjk>
	0x8BB1: '恭' // U+606D <cjk>
	0x8BB2: '挟' // U+631F <cjk>
	0x8BB3: '教' // U+6559 <cjk>
	0x8BB4: '橋' // U+6A4B <cjk>
	0x8BB5: '況' // U+6CC1 <cjk>
	0x8BB6: '狂' // U+72C2 <cjk>
	0x8BB7: '狭' // U+72ED <cjk>
	0x8BB8: '矯' // U+77EF <cjk>
	0x8BB9: '胸' // U+80F8 <cjk>
	0x8BBA: '脅' // U+8105 <cjk>
	0x8BBB: '興' // U+8208 <cjk>
	0x8BBC: '蕎' // U+854E <cjk>
	0x8BBD: '郷' // U+90F7 <cjk>
	0x8BBE: '鏡' // U+93E1 <cjk>
	0x8BBF: '響' // U+97FF <cjk>
	0x8BC0: '饗' // U+9957 <cjk>
	0x8BC1: '驚' // U+9A5A <cjk>
	0x8BC2: '仰' // U+4EF0 <cjk>
	0x8BC3: '凝' // U+51DD <cjk>
	0x8BC4: '尭' // U+5C2D <cjk>
	0x8BC5: '暁' // U+6681 <cjk>
	0x8BC6: '業' // U+696D <cjk>
	0x8BC7: '局' // U+5C40 <cjk>
	0x8BC8: '曲' // U+66F2 <cjk>
	0x8BC9: '極' // U+6975 <cjk>
	0x8BCA: '玉' // U+7389 <cjk>
	0x8BCB: '桐' // U+6850 <cjk>
	0x8BCC: '粁' // U+7C81 <cjk>
	0x8BCD: '僅' // U+50C5 <cjk>
	0x8BCE: '勤' // U+52E4 <cjk>
	0x8BCF: '均' // U+5747 <cjk>
	0x8BD0: '巾' // U+5DFE <cjk>
	0x8BD1: '錦' // U+9326 <cjk>
	0x8BD2: '斤' // U+65A4 <cjk>
	0x8BD3: '欣' // U+6B23 <cjk>
	0x8BD4: '欽' // U+6B3D <cjk>
	0x8BD5: '琴' // U+7434 <cjk>
	0x8BD6: '禁' // U+7981 <cjk>
	0x8BD7: '禽' // U+79BD <cjk>
	0x8BD8: '筋' // U+7B4B <cjk>
	0x8BD9: '緊' // U+7DCA <cjk>
	0x8BDA: '芹' // U+82B9 <cjk>
	0x8BDB: '菌' // U+83CC <cjk>
	0x8BDC: '衿' // U+887F <cjk>
	0x8BDD: '襟' // U+895F <cjk>
	0x8BDE: '謹' // U+8B39 <cjk>
	0x8BDF: '近' // U+8FD1 <cjk>
	0x8BE0: '金' // U+91D1 <cjk>
	0x8BE1: '吟' // U+541F <cjk>
	0x8BE2: '銀' // U+9280 <cjk>
	0x8BE3: '九' // U+4E5D <cjk>
	0x8BE4: '倶' // U+5036 <cjk>
	0x8BE5: '句' // U+53E5 <cjk>
	0x8BE6: '区' // U+533A <cjk>
	0x8BE7: '狗' // U+72D7 <cjk>
	0x8BE8: '玖' // U+7396 <cjk>
	0x8BE9: '矩' // U+77E9 <cjk>
	0x8BEA: '苦' // U+82E6 <cjk>
	0x8BEB: '躯' // U+8EAF <cjk>
	0x8BEC: '駆' // U+99C6 <cjk>
	0x8BED: '駈' // U+99C8 <cjk>
	0x8BEE: '駒' // U+99D2 <cjk>
	0x8BEF: '具' // U+5177 <cjk>
	0x8BF0: '愚' // U+611A <cjk>
	0x8BF1: '虞' // U+865E <cjk>
	0x8BF2: '喰' // U+55B0 <cjk>
	0x8BF3: '空' // U+7A7A <cjk>
	0x8BF4: '偶' // U+5076 <cjk>
	0x8BF5: '寓' // U+5BD3 <cjk>
	0x8BF6: '遇' // U+9047 <cjk>
	0x8BF7: '隅' // U+9685 <cjk>
	0x8BF8: '串' // U+4E32 <cjk>
	0x8BF9: '櫛' // U+6ADB <cjk>
	0x8BFA: '釧' // U+91E7 <cjk>
	0x8BFB: '屑' // U+5C51 <cjk>
	0x8BFC: '屈' // U+5C48 <cjk>
	0x8C40: '掘' // U+6398 <cjk>
	0x8C41: '窟' // U+7A9F <cjk>
	0x8C42: '沓' // U+6C93 <cjk>
	0x8C43: '靴' // U+9774 <cjk>
	0x8C44: '轡' // U+8F61 <cjk>
	0x8C45: '窪' // U+7AAA <cjk>
	0x8C46: '熊' // U+718A <cjk>
	0x8C47: '隈' // U+9688 <cjk>
	0x8C48: '粂' // U+7C82 <cjk>
	0x8C49: '栗' // U+6817 <cjk>
	0x8C4A: '繰' // U+7E70 <cjk>
	0x8C4B: '桑' // U+6851 <cjk>
	0x8C4C: '鍬' // U+936C <cjk>
	0x8C4D: '勲' // U+52F2 <cjk>
	0x8C4E: '君' // U+541B <cjk>
	0x8C4F: '薫' // U+85AB <cjk>
	0x8C50: '訓' // U+8A13 <cjk>
	0x8C51: '群' // U+7FA4 <cjk>
	0x8C52: '軍' // U+8ECD <cjk>
	0x8C53: '郡' // U+90E1 <cjk>
	0x8C54: '卦' // U+5366 <cjk>
	0x8C55: '袈' // U+8888 <cjk>
	0x8C56: '祁' // U+7941 <cjk>
	0x8C57: '係' // U+4FC2 <cjk>
	0x8C58: '傾' // U+50BE <cjk>
	0x8C59: '刑' // U+5211 <cjk>
	0x8C5A: '兄' // U+5144 <cjk>
	0x8C5B: '啓' // U+5553 <cjk>
	0x8C5C: '圭' // U+572D <cjk>
	0x8C5D: '珪' // U+73EA <cjk>
	0x8C5E: '型' // U+578B <cjk>
	0x8C5F: '契' // U+5951 <cjk>
	0x8C60: '形' // U+5F62 <cjk>
	0x8C61: '径' // U+5F84 <cjk>
	0x8C62: '恵' // U+6075 <cjk>
	0x8C63: '慶' // U+6176 <cjk>
	0x8C64: '慧' // U+6167 <cjk>
	0x8C65: '憩' // U+61A9 <cjk>
	0x8C66: '掲' // U+63B2 <cjk>
	0x8C67: '携' // U+643A <cjk>
	0x8C68: '敬' // U+656C <cjk>
	0x8C69: '景' // U+666F <cjk>
	0x8C6A: '桂' // U+6842 <cjk>
	0x8C6B: '渓' // U+6E13 <cjk>
	0x8C6C: '畦' // U+7566 <cjk>
	0x8C6D: '稽' // U+7A3D <cjk>
	0x8C6E: '系' // U+7CFB <cjk>
	0x8C6F: '経' // U+7D4C <cjk>
	0x8C70: '継' // U+7D99 <cjk>
	0x8C71: '繋' // U+7E4B <cjk>
	0x8C72: '罫' // U+7F6B <cjk>
	0x8C73: '茎' // U+830E <cjk>
	0x8C74: '荊' // U+834A <cjk>
	0x8C75: '蛍' // U+86CD <cjk>
	0x8C76: '計' // U+8A08 <cjk>
	0x8C77: '詣' // U+8A63 <cjk>
	0x8C78: '警' // U+8B66 <cjk>
	0x8C79: '軽' // U+8EFD <cjk>
	0x8C7A: '頚' // U+981A <cjk>
	0x8C7B: '鶏' // U+9D8F <cjk>
	0x8C7C: '芸' // U+82B8 <cjk>
	0x8C7D: '迎' // U+8FCE <cjk>
	0x8C7E: '鯨' // U+9BE8 <cjk>
	0x8C80: '劇' // U+5287 <cjk>
	0x8C81: '戟' // U+621F <cjk>
	0x8C82: '撃' // U+6483 <cjk>
	0x8C83: '激' // U+6FC0 <cjk>
	0x8C84: '隙' // U+9699 <cjk>
	0x8C85: '桁' // U+6841 <cjk>
	0x8C86: '傑' // U+5091 <cjk>
	0x8C87: '欠' // U+6B20 <cjk>
	0x8C88: '決' // U+6C7A <cjk>
	0x8C89: '潔' // U+6F54 <cjk>
	0x8C8A: '穴' // U+7A74 <cjk>
	0x8C8B: '結' // U+7D50 <cjk>
	0x8C8C: '血' // U+8840 <cjk>
	0x8C8D: '訣' // U+8A23 <cjk>
	0x8C8E: '月' // U+6708 <cjk>
	0x8C8F: '件' // U+4EF6 <cjk>
	0x8C90: '倹' // U+5039 <cjk>
	0x8C91: '倦' // U+5026 <cjk>
	0x8C92: '健' // U+5065 <cjk>
	0x8C93: '兼' // U+517C <cjk>
	0x8C94: '券' // U+5238 <cjk>
	0x8C95: '剣' // U+5263 <cjk>
	0x8C96: '喧' // U+55A7 <cjk>
	0x8C97: '圏' // U+570F <cjk>
	0x8C98: '堅' // U+5805 <cjk>
	0x8C99: '嫌' // U+5ACC <cjk>
	0x8C9A: '建' // U+5EFA <cjk>
	0x8C9B: '憲' // U+61B2 <cjk>
	0x8C9C: '懸' // U+61F8 <cjk>
	0x8C9D: '拳' // U+62F3 <cjk>
	0x8C9E: '捲' // U+6372 <cjk>
	0x8C9F: '検' // U+691C <cjk>
	0x8CA0: '権' // U+6A29 <cjk>
	0x8CA1: '牽' // U+727D <cjk>
	0x8CA2: '犬' // U+72AC <cjk>
	0x8CA3: '献' // U+732E <cjk>
	0x8CA4: '研' // U+7814 <cjk>
	0x8CA5: '硯' // U+786F <cjk>
	0x8CA6: '絹' // U+7D79 <cjk>
	0x8CA7: '県' // U+770C <cjk>
	0x8CA8: '肩' // U+80A9 <cjk>
	0x8CA9: '見' // U+898B <cjk>
	0x8CAA: '謙' // U+8B19 <cjk>
	0x8CAB: '賢' // U+8CE2 <cjk>
	0x8CAC: '軒' // U+8ED2 <cjk>
	0x8CAD: '遣' // U+9063 <cjk>
	0x8CAE: '鍵' // U+9375 <cjk>
	0x8CAF: '険' // U+967A <cjk>
	0x8CB0: '顕' // U+9855 <cjk>
	0x8CB1: '験' // U+9A13 <cjk>
	0x8CB2: '鹸' // U+9E78 <cjk>
	0x8CB3: '元' // U+5143 <cjk>
	0x8CB4: '原' // U+539F <cjk>
	0x8CB5: '厳' // U+53B3 <cjk>
	0x8CB6: '幻' // U+5E7B <cjk>
	0x8CB7: '弦' // U+5F26 <cjk>
	0x8CB8: '減' // U+6E1B <cjk>
	0x8CB9: '源' // U+6E90 <cjk>
	0x8CBA: '玄' // U+7384 <cjk>
	0x8CBB: '現' // U+73FE <cjk>
	0x8CBC: '絃' // U+7D43 <cjk>
	0x8CBD: '舷' // U+8237 <cjk>
	0x8CBE: '言' // U+8A00 <cjk>
	0x8CBF: '諺' // U+8AFA <cjk>
	0x8CC0: '限' // U+9650 <cjk>
	0x8CC1: '乎' // U+4E4E <cjk>
	0x8CC2: '個' // U+500B <cjk>
	0x8CC3: '古' // U+53E4 <cjk>
	0x8CC4: '呼' // U+547C <cjk>
	0x8CC5: '固' // U+56FA <cjk>
	0x8CC6: '姑' // U+59D1 <cjk>
	0x8CC7: '孤' // U+5B64 <cjk>
	0x8CC8: '己' // U+5DF1 <cjk>
	0x8CC9: '庫' // U+5EAB <cjk>
	0x8CCA: '弧' // U+5F27 <cjk>
	0x8CCB: '戸' // U+6238 <cjk>
	0x8CCC: '故' // U+6545 <cjk>
	0x8CCD: '枯' // U+67AF <cjk>
	0x8CCE: '湖' // U+6E56 <cjk>
	0x8CCF: '狐' // U+72D0 <cjk>
	0x8CD0: '糊' // U+7CCA <cjk>
	0x8CD1: '袴' // U+88B4 <cjk>
	0x8CD2: '股' // U+80A1 <cjk>
	0x8CD3: '胡' // U+80E1 <cjk>
	0x8CD4: '菰' // U+83F0 <cjk>
	0x8CD5: '虎' // U+864E <cjk>
	0x8CD6: '誇' // U+8A87 <cjk>
	0x8CD7: '跨' // U+8DE8 <cjk>
	0x8CD8: '鈷' // U+9237 <cjk>
	0x8CD9: '雇' // U+96C7 <cjk>
	0x8CDA: '顧' // U+9867 <cjk>
	0x8CDB: '鼓' // U+9F13 <cjk>
	0x8CDC: '五' // U+4E94 <cjk>
	0x8CDD: '互' // U+4E92 <cjk>
	0x8CDE: '伍' // U+4F0D <cjk>
	0x8CDF: '午' // U+5348 <cjk>
	0x8CE0: '呉' // U+5449 <cjk>
	0x8CE1: '吾' // U+543E <cjk>
	0x8CE2: '娯' // U+5A2F <cjk>
	0x8CE3: '後' // U+5F8C <cjk>
	0x8CE4: '御' // U+5FA1 <cjk>
	0x8CE5: '悟' // U+609F <cjk>
	0x8CE6: '梧' // U+68A7 <cjk>
	0x8CE7: '檎' // U+6A8E <cjk>
	0x8CE8: '瑚' // U+745A <cjk>
	0x8CE9: '碁' // U+7881 <cjk>
	0x8CEA: '語' // U+8A9E <cjk>
	0x8CEB: '誤' // U+8AA4 <cjk>
	0x8CEC: '護' // U+8B77 <cjk>
	0x8CED: '醐' // U+9190 <cjk>
	0x8CEE: '乞' // U+4E5E <cjk>
	0x8CEF: '鯉' // U+9BC9 <cjk>
	0x8CF0: '交' // U+4EA4 <cjk>
	0x8CF1: '佼' // U+4F7C <cjk>
	0x8CF2: '侯' // U+4FAF <cjk>
	0x8CF3: '候' // U+5019 <cjk>
	0x8CF4: '倖' // U+5016 <cjk>
	0x8CF5: '光' // U+5149 <cjk>
	0x8CF6: '公' // U+516C <cjk>
	0x8CF7: '功' // U+529F <cjk>
	0x8CF8: '効' // U+52B9 <cjk>
	0x8CF9: '勾' // U+52FE <cjk>
	0x8CFA: '厚' // U+539A <cjk>
	0x8CFB: '口' // U+53E3 <cjk>
	0x8CFC: '向' // U+5411 <cjk>
	0x8D40: '后' // U+540E <cjk>
	0x8D41: '喉' // U+5589 <cjk>
	0x8D42: '坑' // U+5751 <cjk>
	0x8D43: '垢' // U+57A2 <cjk>
	0x8D44: '好' // U+597D <cjk>
	0x8D45: '孔' // U+5B54 <cjk>
	0x8D46: '孝' // U+5B5D <cjk>
	0x8D47: '宏' // U+5B8F <cjk>
	0x8D48: '工' // U+5DE5 <cjk>
	0x8D49: '巧' // U+5DE7 <cjk>
	0x8D4A: '巷' // U+5DF7 <cjk>
	0x8D4B: '幸' // U+5E78 <cjk>
	0x8D4C: '広' // U+5E83 <cjk>
	0x8D4D: '庚' // U+5E9A <cjk>
	0x8D4E: '康' // U+5EB7 <cjk>
	0x8D4F: '弘' // U+5F18 <cjk>
	0x8D50: '恒' // U+6052 <cjk>
	0x8D51: '慌' // U+614C <cjk>
	0x8D52: '抗' // U+6297 <cjk>
	0x8D53: '拘' // U+62D8 <cjk>
	0x8D54: '控' // U+63A7 <cjk>
	0x8D55: '攻' // U+653B <cjk>
	0x8D56: '昂' // U+6602 <cjk>
	0x8D57: '晃' // U+6643 <cjk>
	0x8D58: '更' // U+66F4 <cjk>
	0x8D59: '杭' // U+676D <cjk>
	0x8D5A: '校' // U+6821 <cjk>
	0x8D5B: '梗' // U+6897 <cjk>
	0x8D5C: '構' // U+69CB <cjk>
	0x8D5D: '江' // U+6C5F <cjk>
	0x8D5E: '洪' // U+6D2A <cjk>
	0x8D5F: '浩' // U+6D69 <cjk>
	0x8D60: '港' // U+6E2F <cjk>
	0x8D61: '溝' // U+6E9D <cjk>
	0x8D62: '甲' // U+7532 <cjk>
	0x8D63: '皇' // U+7687 <cjk>
	0x8D64: '硬' // U+786C <cjk>
	0x8D65: '稿' // U+7A3F <cjk>
	0x8D66: '糠' // U+7CE0 <cjk>
	0x8D67: '紅' // U+7D05 <cjk>
	0x8D68: '紘' // U+7D18 <cjk>
	0x8D69: '絞' // U+7D5E <cjk>
	0x8D6A: '綱' // U+7DB1 <cjk>
	0x8D6B: '耕' // U+8015 <cjk>
	0x8D6C: '考' // U+8003 <cjk>
	0x8D6D: '肯' // U+80AF <cjk>
	0x8D6E: '肱' // U+80B1 <cjk>
	0x8D6F: '腔' // U+8154 <cjk>
	0x8D70: '膏' // U+818F <cjk>
	0x8D71: '航' // U+822A <cjk>
	0x8D72: '荒' // U+8352 <cjk>
	0x8D73: '行' // U+884C <cjk>
	0x8D74: '衡' // U+8861 <cjk>
	0x8D75: '講' // U+8B1B <cjk>
	0x8D76: '貢' // U+8CA2 <cjk>
	0x8D77: '購' // U+8CFC <cjk>
	0x8D78: '郊' // U+90CA <cjk>
	0x8D79: '酵' // U+9175 <cjk>
	0x8D7A: '鉱' // U+9271 <cjk>
	0x8D7B: '砿' // U+783F <cjk>
	0x8D7C: '鋼' // U+92FC <cjk>
	0x8D7D: '閤' // U+95A4 <cjk>
	0x8D7E: '降' // U+964D <cjk>
	0x8D80: '項' // U+9805 <cjk>
	0x8D81: '香' // U+9999 <cjk>
	0x8D82: '高' // U+9AD8 <cjk>
	0x8D83: '鴻' // U+9D3B <cjk>
	0x8D84: '剛' // U+525B <cjk>
	0x8D85: '劫' // U+52AB <cjk>
	0x8D86: '号' // U+53F7 <cjk>
	0x8D87: '合' // U+5408 <cjk>
	0x8D88: '壕' // U+58D5 <cjk>
	0x8D89: '拷' // U+62F7 <cjk>
	0x8D8A: '濠' // U+6FE0 <cjk>
	0x8D8B: '豪' // U+8C6A <cjk>
	0x8D8C: '轟' // U+8F5F <cjk>
	0x8D8D: '麹' // U+9EB9 <cjk>
	0x8D8E: '克' // U+514B <cjk>
	0x8D8F: '刻' // U+523B <cjk>
	0x8D90: '告' // U+544A <cjk>
	0x8D91: '国' // U+56FD <cjk>
	0x8D92: '穀' // U+7A40 <cjk>
	0x8D93: '酷' // U+9177 <cjk>
	0x8D94: '鵠' // U+9D60 <cjk>
	0x8D95: '黒' // U+9ED2 <cjk>
	0x8D96: '獄' // U+7344 <cjk>
	0x8D97: '漉' // U+6F09 <cjk>
	0x8D98: '腰' // U+8170 <cjk>
	0x8D99: '甑' // U+7511 <cjk>
	0x8D9A: '忽' // U+5FFD <cjk>
	0x8D9B: '惚' // U+60DA <cjk>
	0x8D9C: '骨' // U+9AA8 <cjk>
	0x8D9D: '狛' // U+72DB <cjk>
	0x8D9E: '込' // U+8FBC <cjk>
	0x8D9F: '此' // U+6B64 <cjk>
	0x8DA0: '頃' // U+9803 <cjk>
	0x8DA1: '今' // U+4ECA <cjk>
	0x8DA2: '困' // U+56F0 <cjk>
	0x8DA3: '坤' // U+5764 <cjk>
	0x8DA4: '墾' // U+58BE <cjk>
	0x8DA5: '婚' // U+5A5A <cjk>
	0x8DA6: '恨' // U+6068 <cjk>
	0x8DA7: '懇' // U+61C7 <cjk>
	0x8DA8: '昏' // U+660F <cjk>
	0x8DA9: '昆' // U+6606 <cjk>
	0x8DAA: '根' // U+6839 <cjk>
	0x8DAB: '梱' // U+68B1 <cjk>
	0x8DAC: '混' // U+6DF7 <cjk>
	0x8DAD: '痕' // U+75D5 <cjk>
	0x8DAE: '紺' // U+7D3A <cjk>
	0x8DAF: '艮' // U+826E <cjk>
	0x8DB0: '魂' // U+9B42 <cjk>
	0x8DB1: '些' // U+4E9B <cjk>
	0x8DB2: '佐' // U+4F50 <cjk>
	0x8DB3: '叉' // U+53C9 <cjk>
	0x8DB4: '唆' // U+5506 <cjk>
	0x8DB5: '嵯' // U+5D6F <cjk>
	0x8DB6: '左' // U+5DE6 <cjk>
	0x8DB7: '差' // U+5DEE <cjk>
	0x8DB8: '査' // U+67FB <cjk>
	0x8DB9: '沙' // U+6C99 <cjk>
	0x8DBA: '瑳' // U+7473 <cjk>
	0x8DBB: '砂' // U+7802 <cjk>
	0x8DBC: '詐' // U+8A50 <cjk>
	0x8DBD: '鎖' // U+9396 <cjk>
	0x8DBE: '裟' // U+88DF <cjk>
	0x8DBF: '坐' // U+5750 <cjk>
	0x8DC0: '座' // U+5EA7 <cjk>
	0x8DC1: '挫' // U+632B <cjk>
	0x8DC2: '債' // U+50B5 <cjk>
	0x8DC3: '催' // U+50AC <cjk>
	0x8DC4: '再' // U+518D <cjk>
	0x8DC5: '最' // U+6700 <cjk>
	0x8DC6: '哉' // U+54C9 <cjk>
	0x8DC7: '塞' // U+585E <cjk>
	0x8DC8: '妻' // U+59BB <cjk>
	0x8DC9: '宰' // U+5BB0 <cjk>
	0x8DCA: '彩' // U+5F69 <cjk>
	0x8DCB: '才' // U+624D <cjk>
	0x8DCC: '採' // U+63A1 <cjk>
	0x8DCD: '栽' // U+683D <cjk>
	0x8DCE: '歳' // U+6B73 <cjk>
	0x8DCF: '済' // U+6E08 <cjk>
	0x8DD0: '災' // U+707D <cjk>
	0x8DD1: '采' // U+91C7 <cjk>
	0x8DD2: '犀' // U+7280 <cjk>
	0x8DD3: '砕' // U+7815 <cjk>
	0x8DD4: '砦' // U+7826 <cjk>
	0x8DD5: '祭' // U+796D <cjk>
	0x8DD6: '斎' // U+658E <cjk>
	0x8DD7: '細' // U+7D30 <cjk>
	0x8DD8: '菜' // U+83DC <cjk>
	0x8DD9: '裁' // U+88C1 <cjk>
	0x8DDA: '載' // U+8F09 <cjk>
	0x8DDB: '際' // U+969B <cjk>
	0x8DDC: '剤' // U+5264 <cjk>
	0x8DDD: '在' // U+5728 <cjk>
	0x8DDE: '材' // U+6750 <cjk>
	0x8DDF: '罪' // U+7F6A <cjk>
	0x8DE0: '財' // U+8CA1 <cjk>
	0x8DE1: '冴' // U+51B4 <cjk>
	0x8DE2: '坂' // U+5742 <cjk>
	0x8DE3: '阪' // U+962A <cjk>
	0x8DE4: '堺' // U+583A <cjk>
	0x8DE5: '榊' // U+698A <cjk>
	0x8DE6: '肴' // U+80B4 <cjk>
	0x8DE7: '咲' // U+54B2 <cjk>
	0x8DE8: '崎' // U+5D0E <cjk>
	0x8DE9: '埼' // U+57FC <cjk>
	0x8DEA: '碕' // U+7895 <cjk>
	0x8DEB: '鷺' // U+9DFA <cjk>
	0x8DEC: '作' // U+4F5C <cjk>
	0x8DED: '削' // U+524A <cjk>
	0x8DEE: '咋' // U+548B <cjk>
	0x8DEF: '搾' // U+643E <cjk>
	0x8DF0: '昨' // U+6628 <cjk>
	0x8DF1: '朔' // U+6714 <cjk>
	0x8DF2: '柵' // U+67F5 <cjk>
	0x8DF3: '窄' // U+7A84 <cjk>
	0x8DF4: '策' // U+7B56 <cjk>
	0x8DF5: '索' // U+7D22 <cjk>
	0x8DF6: '錯' // U+932F <cjk>
	0x8DF7: '桜' // U+685C <cjk>
	0x8DF8: '鮭' // U+9BAD <cjk>
	0x8DF9: '笹' // U+7B39 <cjk>
	0x8DFA: '匙' // U+5319 <cjk>
	0x8DFB: '冊' // U+518A <cjk>
	0x8DFC: '刷' // U+5237 <cjk>
	0x8E40: '察' // U+5BDF <cjk>
	0x8E41: '拶' // U+62F6 <cjk>
	0x8E42: '撮' // U+64AE <cjk>
	0x8E43: '擦' // U+64E6 <cjk>
	0x8E44: '札' // U+672D <cjk>
	0x8E45: '殺' // U+6BBA <cjk>
	0x8E46: '薩' // U+85A9 <cjk>
	0x8E47: '雑' // U+96D1 <cjk>
	0x8E48: '皐' // U+7690 <cjk>
	0x8E49: '鯖' // U+9BD6 <cjk>
	0x8E4A: '捌' // U+634C <cjk>
	0x8E4B: '錆' // U+9306 <cjk>
	0x8E4C: '鮫' // U+9BAB <cjk>
	0x8E4D: '皿' // U+76BF <cjk>
	0x8E4E: '晒' // U+6652 <cjk>
	0x8E4F: '三' // U+4E09 <cjk>
	0x8E50: '傘' // U+5098 <cjk>
	0x8E51: '参' // U+53C2 <cjk>
	0x8E52: '山' // U+5C71 <cjk>
	0x8E53: '惨' // U+60E8 <cjk>
	0x8E54: '撒' // U+6492 <cjk>
	0x8E55: '散' // U+6563 <cjk>
	0x8E56: '桟' // U+685F <cjk>
	0x8E57: '燦' // U+71E6 <cjk>
	0x8E58: '珊' // U+73CA <cjk>
	0x8E59: '産' // U+7523 <cjk>
	0x8E5A: '算' // U+7B97 <cjk>
	0x8E5B: '纂' // U+7E82 <cjk>
	0x8E5C: '蚕' // U+8695 <cjk>
	0x8E5D: '讃' // U+8B83 <cjk>
	0x8E5E: '賛' // U+8CDB <cjk>
	0x8E5F: '酸' // U+9178 <cjk>
	0x8E60: '餐' // U+9910 <cjk>
	0x8E61: '斬' // U+65AC <cjk>
	0x8E62: '暫' // U+66AB <cjk>
	0x8E63: '残' // U+6B8B <cjk>
	0x8E64: '仕' // U+4ED5 <cjk>
	0x8E65: '仔' // U+4ED4 <cjk>
	0x8E66: '伺' // U+4F3A <cjk>
	0x8E67: '使' // U+4F7F <cjk>
	0x8E68: '刺' // U+523A <cjk>
	0x8E69: '司' // U+53F8 <cjk>
	0x8E6A: '史' // U+53F2 <cjk>
	0x8E6B: '嗣' // U+55E3 <cjk>
	0x8E6C: '四' // U+56DB <cjk>
	0x8E6D: '士' // U+58EB <cjk>
	0x8E6E: '始' // U+59CB <cjk>
	0x8E6F: '姉' // U+59C9 <cjk>
	0x8E70: '姿' // U+59FF <cjk>
	0x8E71: '子' // U+5B50 <cjk>
	0x8E72: '屍' // U+5C4D <cjk>
	0x8E73: '市' // U+5E02 <cjk>
	0x8E74: '師' // U+5E2B <cjk>
	0x8E75: '志' // U+5FD7 <cjk>
	0x8E76: '思' // U+601D <cjk>
	0x8E77: '指' // U+6307 <cjk>
	0x8E78: '支' // U+652F <cjk>
	0x8E79: '孜' // U+5B5C <cjk>
	0x8E7A: '斯' // U+65AF <cjk>
	0x8E7B: '施' // U+65BD <cjk>
	0x8E7C: '旨' // U+65E8 <cjk>
	0x8E7D: '枝' // U+679D <cjk>
	0x8E7E: '止' // U+6B62 <cjk>
	0x8E80: '死' // U+6B7B <cjk>
	0x8E81: '氏' // U+6C0F <cjk>
	0x8E82: '獅' // U+7345 <cjk>
	0x8E83: '祉' // U+7949 <cjk>
	0x8E84: '私' // U+79C1 <cjk>
	0x8E85: '糸' // U+7CF8 <cjk>
	0x8E86: '紙' // U+7D19 <cjk>
	0x8E87: '紫' // U+7D2B <cjk>
	0x8E88: '肢' // U+80A2 <cjk>
	0x8E89: '脂' // U+8102 <cjk>
	0x8E8A: '至' // U+81F3 <cjk>
	0x8E8B: '視' // U+8996 <cjk>
	0x8E8C: '詞' // U+8A5E <cjk>
	0x8E8D: '詩' // U+8A69 <cjk>
	0x8E8E: '試' // U+8A66 <cjk>
	0x8E8F: '誌' // U+8A8C <cjk>
	0x8E90: '諮' // U+8AEE <cjk>
	0x8E91: '資' // U+8CC7 <cjk>
	0x8E92: '賜' // U+8CDC <cjk>
	0x8E93: '雌' // U+96CC <cjk>
	0x8E94: '飼' // U+98FC <cjk>
	0x8E95: '歯' // U+6B6F <cjk>
	0x8E96: '事' // U+4E8B <cjk>
	0x8E97: '似' // U+4F3C <cjk>
	0x8E98: '侍' // U+4F8D <cjk>
	0x8E99: '児' // U+5150 <cjk>
	0x8E9A: '字' // U+5B57 <cjk>
	0x8E9B: '寺' // U+5BFA <cjk>
	0x8E9C: '慈' // U+6148 <cjk>
	0x8E9D: '持' // U+6301 <cjk>
	0x8E9E: '時' // U+6642 <cjk>
	0x8E9F: '次' // U+6B21 <cjk>
	0x8EA0: '滋' // U+6ECB <cjk>
	0x8EA1: '治' // U+6CBB <cjk>
	0x8EA2: '爾' // U+723E <cjk>
	0x8EA3: '璽' // U+74BD <cjk>
	0x8EA4: '痔' // U+75D4 <cjk>
	0x8EA5: '磁' // U+78C1 <cjk>
	0x8EA6: '示' // U+793A <cjk>
	0x8EA7: '而' // U+800C <cjk>
	0x8EA8: '耳' // U+8033 <cjk>
	0x8EA9: '自' // U+81EA <cjk>
	0x8EAA: '蒔' // U+8494 <cjk>
	0x8EAB: '辞' // U+8F9E <cjk>
	0x8EAC: '汐' // U+6C50 <cjk>
	0x8EAD: '鹿' // U+9E7F <cjk>
	0x8EAE: '式' // U+5F0F <cjk>
	0x8EAF: '識' // U+8B58 <cjk>
	0x8EB0: '鴫' // U+9D2B <cjk>
	0x8EB1: '竺' // U+7AFA <cjk>
	0x8EB2: '軸' // U+8EF8 <cjk>
	0x8EB3: '宍' // U+5B8D <cjk>
	0x8EB4: '雫' // U+96EB <cjk>
	0x8EB5: '七' // U+4E03 <cjk>
	0x8EB6: '叱' // U+53F1 <cjk>
	0x8EB7: '執' // U+57F7 <cjk>
	0x8EB8: '失' // U+5931 <cjk>
	0x8EB9: '嫉' // U+5AC9 <cjk>
	0x8EBA: '室' // U+5BA4 <cjk>
	0x8EBB: '悉' // U+6089 <cjk>
	0x8EBC: '湿' // U+6E7F <cjk>
	0x8EBD: '漆' // U+6F06 <cjk>
	0x8EBE: '疾' // U+75BE <cjk>
	0x8EBF: '質' // U+8CEA <cjk>
	0x8EC0: '実' // U+5B9F <cjk>
	0x8EC1: '蔀' // U+8500 <cjk>
	0x8EC2: '篠' // U+7BE0 <cjk>
	0x8EC3: '偲' // U+5072 <cjk>
	0x8EC4: '柴' // U+67F4 <cjk>
	0x8EC5: '芝' // U+829D <cjk>
	0x8EC6: '屡' // U+5C61 <cjk>
	0x8EC7: '蕊' // U+854A <cjk>
	0x8EC8: '縞' // U+7E1E <cjk>
	0x8EC9: '舎' // U+820E <cjk>
	0x8ECA: '写' // U+5199 <cjk>
	0x8ECB: '射' // U+5C04 <cjk>
	0x8ECC: '捨' // U+6368 <cjk>
	0x8ECD: '赦' // U+8D66 <cjk>
	0x8ECE: '斜' // U+659C <cjk>
	0x8ECF: '煮' // U+716E <cjk>
	0x8ED0: '社' // U+793E <cjk>
	0x8ED1: '紗' // U+7D17 <cjk>
	0x8ED2: '者' // U+8005 <cjk>
	0x8ED3: '謝' // U+8B1D <cjk>
	0x8ED4: '車' // U+8ECA <cjk>
	0x8ED5: '遮' // U+906E <cjk>
	0x8ED6: '蛇' // U+86C7 <cjk>
	0x8ED7: '邪' // U+90AA <cjk>
	0x8ED8: '借' // U+501F <cjk>
	0x8ED9: '勺' // U+52FA <cjk>
	0x8EDA: '尺' // U+5C3A <cjk>
	0x8EDB: '杓' // U+6753 <cjk>
	0x8EDC: '灼' // U+707C <cjk>
	0x8EDD: '爵' // U+7235 <cjk>
	0x8EDE: '酌' // U+914C <cjk>
	0x8EDF: '釈' // U+91C8 <cjk>
	0x8EE0: '錫' // U+932B <cjk>
	0x8EE1: '若' // U+82E5 <cjk>
	0x8EE2: '寂' // U+5BC2 <cjk>
	0x8EE3: '弱' // U+5F31 <cjk>
	0x8EE4: '惹' // U+60F9 <cjk>
	0x8EE5: '主' // U+4E3B <cjk>
	0x8EE6: '取' // U+53D6 <cjk>
	0x8EE7: '守' // U+5B88 <cjk>
	0x8EE8: '手' // U+624B <cjk>
	0x8EE9: '朱' // U+6731 <cjk>
	0x8EEA: '殊' // U+6B8A <cjk>
	0x8EEB: '狩' // U+72E9 <cjk>
	0x8EEC: '珠' // U+73E0 <cjk>
	0x8EED: '種' // U+7A2E <cjk>
	0x8EEE: '腫' // U+816B <cjk>
	0x8EEF: '趣' // U+8DA3 <cjk>
	0x8EF0: '酒' // U+9152 <cjk>
	0x8EF1: '首' // U+9996 <cjk>
	0x8EF2: '儒' // U+5112 <cjk>
	0x8EF3: '受' // U+53D7 <cjk>
	0x8EF4: '呪' // U+546A <cjk>
	0x8EF5: '寿' // U+5BFF <cjk>
	0x8EF6: '授' // U+6388 <cjk>
	0x8EF7: '樹' // U+6A39 <cjk>
	0x8EF8: '綬' // U+7DAC <cjk>
	0x8EF9: '需' // U+9700 <cjk>
	0x8EFA: '囚' // U+56DA <cjk>
	0x8EFB: '収' // U+53CE <cjk>
	0x8EFC: '周' // U+5468 <cjk>
	0x8F40: '宗' // U+5B97 <cjk>
	0x8F41: '就' // U+5C31 <cjk>
	0x8F42: '州' // U+5DDE <cjk>
	0x8F43: '修' // U+4FEE <cjk>
	0x8F44: '愁' // U+6101 <cjk>
	0x8F45: '拾' // U+62FE <cjk>
	0x8F46: '洲' // U+6D32 <cjk>
	0x8F47: '秀' // U+79C0 <cjk>
	0x8F48: '秋' // U+79CB <cjk>
	0x8F49: '終' // U+7D42 <cjk>
	0x8F4A: '繍' // U+7E4D <cjk>
	0x8F4B: '習' // U+7FD2 <cjk>
	0x8F4C: '臭' // U+81ED <cjk>
	0x8F4D: '舟' // U+821F <cjk>
	0x8F4E: '蒐' // U+8490 <cjk>
	0x8F4F: '衆' // U+8846 <cjk>
	0x8F50: '襲' // U+8972 <cjk>
	0x8F51: '讐' // U+8B90 <cjk>
	0x8F52: '蹴' // U+8E74 <cjk>
	0x8F53: '輯' // U+8F2F <cjk>
	0x8F54: '週' // U+9031 <cjk>
	0x8F55: '酋' // U+914B <cjk>
	0x8F56: '酬' // U+916C <cjk>
	0x8F57: '集' // U+96C6 <cjk>
	0x8F58: '醜' // U+919C <cjk>
	0x8F59: '什' // U+4EC0 <cjk>
	0x8F5A: '住' // U+4F4F <cjk>
	0x8F5B: '充' // U+5145 <cjk>
	0x8F5C: '十' // U+5341 <cjk>
	0x8F5D: '従' // U+5F93 <cjk>
	0x8F5E: '戎' // U+620E <cjk>
	0x8F5F: '柔' // U+67D4 <cjk>
	0x8F60: '汁' // U+6C41 <cjk>
	0x8F61: '渋' // U+6E0B <cjk>
	0x8F62: '獣' // U+7363 <cjk>
	0x8F63: '縦' // U+7E26 <cjk>
	0x8F64: '重' // U+91CD <cjk>
	0x8F65: '銃' // U+9283 <cjk>
	0x8F66: '叔' // U+53D4 <cjk>
	0x8F67: '夙' // U+5919 <cjk>
	0x8F68: '宿' // U+5BBF <cjk>
	0x8F69: '淑' // U+6DD1 <cjk>
	0x8F6A: '祝' // U+795D <cjk>
	0x8F6B: '縮' // U+7E2E <cjk>
	0x8F6C: '粛' // U+7C9B <cjk>
	0x8F6D: '塾' // U+587E <cjk>
	0x8F6E: '熟' // U+719F <cjk>
	0x8F6F: '出' // U+51FA <cjk>
	0x8F70: '術' // U+8853 <cjk>
	0x8F71: '述' // U+8FF0 <cjk>
	0x8F72: '俊' // U+4FCA <cjk>
	0x8F73: '峻' // U+5CFB <cjk>
	0x8F74: '春' // U+6625 <cjk>
	0x8F75: '瞬' // U+77AC <cjk>
	0x8F76: '竣' // U+7AE3 <cjk>
	0x8F77: '舜' // U+821C <cjk>
	0x8F78: '駿' // U+99FF <cjk>
	0x8F79: '准' // U+51C6 <cjk>
	0x8F7A: '循' // U+5FAA <cjk>
	0x8F7B: '旬' // U+65EC <cjk>
	0x8F7C: '楯' // U+696F <cjk>
	0x8F7D: '殉' // U+6B89 <cjk>
	0x8F7E: '淳' // U+6DF3 <cjk>
	0x8F80: '準' // U+6E96 <cjk>
	0x8F81: '潤' // U+6F64 <cjk>
	0x8F82: '盾' // U+76FE <cjk>
	0x8F83: '純' // U+7D14 <cjk>
	0x8F84: '巡' // U+5DE1 <cjk>
	0x8F85: '遵' // U+9075 <cjk>
	0x8F86: '醇' // U+9187 <cjk>
	0x8F87: '順' // U+9806 <cjk>
	0x8F88: '処' // U+51E6 <cjk>
	0x8F89: '初' // U+521D <cjk>
	0x8F8A: '所' // U+6240 <cjk>
	0x8F8B: '暑' // U+6691 <cjk>
	0x8F8C: '曙' // U+66D9 <cjk>
	0x8F8D: '渚' // U+6E1A <cjk>
	0x8F8E: '庶' // U+5EB6 <cjk>
	0x8F8F: '緒' // U+7DD2 <cjk>
	0x8F90: '署' // U+7F72 <cjk>
	0x8F91: '書' // U+66F8 <cjk>
	0x8F92: '薯' // U+85AF <cjk>
	0x8F93: '藷' // U+85F7 <cjk>
	0x8F94: '諸' // U+8AF8 <cjk>
	0x8F95: '助' // U+52A9 <cjk>
	0x8F96: '叙' // U+53D9 <cjk>
	0x8F97: '女' // U+5973 <cjk>
	0x8F98: '序' // U+5E8F <cjk>
	0x8F99: '徐' // U+5F90 <cjk>
	0x8F9A: '恕' // U+6055 <cjk>
	0x8F9B: '鋤' // U+92E4 <cjk>
	0x8F9C: '除' // U+9664 <cjk>
	0x8F9D: '傷' // U+50B7 <cjk>
	0x8F9E: '償' // U+511F <cjk>
	0x8F9F: '勝' // U+52DD <cjk>
	0x8FA0: '匠' // U+5320 <cjk>
	0x8FA1: '升' // U+5347 <cjk>
	0x8FA2: '召' // U+53EC <cjk>
	0x8FA3: '哨' // U+54E8 <cjk>
	0x8FA4: '商' // U+5546 <cjk>
	0x8FA5: '唱' // U+5531 <cjk>
	0x8FA6: '嘗' // U+5617 <cjk>
	0x8FA7: '奨' // U+5968 <cjk>
	0x8FA8: '妾' // U+59BE <cjk>
	0x8FA9: '娼' // U+5A3C <cjk>
	0x8FAA: '宵' // U+5BB5 <cjk>
	0x8FAB: '将' // U+5C06 <cjk>
	0x8FAC: '小' // U+5C0F <cjk>
	0x8FAD: '少' // U+5C11 <cjk>
	0x8FAE: '尚' // U+5C1A <cjk>
	0x8FAF: '庄' // U+5E84 <cjk>
	0x8FB0: '床' // U+5E8A <cjk>
	0x8FB1: '廠' // U+5EE0 <cjk>
	0x8FB2: '彰' // U+5F70 <cjk>
	0x8FB3: '承' // U+627F <cjk>
	0x8FB4: '抄' // U+6284 <cjk>
	0x8FB5: '招' // U+62DB <cjk>
	0x8FB6: '掌' // U+638C <cjk>
	0x8FB7: '捷' // U+6377 <cjk>
	0x8FB8: '昇' // U+6607 <cjk>
	0x8FB9: '昌' // U+660C <cjk>
	0x8FBA: '昭' // U+662D <cjk>
	0x8FBB: '晶' // U+6676 <cjk>
	0x8FBC: '松' // U+677E <cjk>
	0x8FBD: '梢' // U+68A2 <cjk>
	0x8FBE: '樟' // U+6A1F <cjk>
	0x8FBF: '樵' // U+6A35 <cjk>
	0x8FC0: '沼' // U+6CBC <cjk>
	0x8FC1: '消' // U+6D88 <cjk>
	0x8FC2: '渉' // U+6E09 <cjk>
	0x8FC3: '湘' // U+6E58 <cjk>
	0x8FC4: '焼' // U+713C <cjk>
	0x8FC5: '焦' // U+7126 <cjk>
	0x8FC6: '照' // U+7167 <cjk>
	0x8FC7: '症' // U+75C7 <cjk>
	0x8FC8: '省' // U+7701 <cjk>
	0x8FC9: '硝' // U+785D <cjk>
	0x8FCA: '礁' // U+7901 <cjk>
	0x8FCB: '祥' // U+7965 <cjk>
	0x8FCC: '称' // U+79F0 <cjk>
	0x8FCD: '章' // U+7AE0 <cjk>
	0x8FCE: '笑' // U+7B11 <cjk>
	0x8FCF: '粧' // U+7CA7 <cjk>
	0x8FD0: '紹' // U+7D39 <cjk>
	0x8FD1: '肖' // U+8096 <cjk>
	0x8FD2: '菖' // U+83D6 <cjk>
	0x8FD3: '蒋' // U+848B <cjk>
	0x8FD4: '蕉' // U+8549 <cjk>
	0x8FD5: '衝' // U+885D <cjk>
	0x8FD6: '裳' // U+88F3 <cjk>
	0x8FD7: '訟' // U+8A1F <cjk>
	0x8FD8: '証' // U+8A3C <cjk>
	0x8FD9: '詔' // U+8A54 <cjk>
	0x8FDA: '詳' // U+8A73 <cjk>
	0x8FDB: '象' // U+8C61 <cjk>
	0x8FDC: '賞' // U+8CDE <cjk>
	0x8FDD: '醤' // U+91A4 <cjk>
	0x8FDE: '鉦' // U+9266 <cjk>
	0x8FDF: '鍾' // U+937E <cjk>
	0x8FE0: '鐘' // U+9418 <cjk>
	0x8FE1: '障' // U+969C <cjk>
	0x8FE2: '鞘' // U+9798 <cjk>
	0x8FE3: '上' // U+4E0A <cjk>
	0x8FE4: '丈' // U+4E08 <cjk>
	0x8FE5: '丞' // U+4E1E <cjk>
	0x8FE6: '乗' // U+4E57 <cjk>
	0x8FE7: '冗' // U+5197 <cjk>
	0x8FE8: '剰' // U+5270 <cjk>
	0x8FE9: '城' // U+57CE <cjk>
	0x8FEA: '場' // U+5834 <cjk>
	0x8FEB: '壌' // U+58CC <cjk>
	0x8FEC: '嬢' // U+5B22 <cjk>
	0x8FED: '常' // U+5E38 <cjk>
	0x8FEE: '情' // U+60C5 <cjk>
	0x8FEF: '擾' // U+64FE <cjk>
	0x8FF0: '条' // U+6761 <cjk>
	0x8FF1: '杖' // U+6756 <cjk>
	0x8FF2: '浄' // U+6D44 <cjk>
	0x8FF3: '状' // U+72B6 <cjk>
	0x8FF4: '畳' // U+7573 <cjk>
	0x8FF5: '穣' // U+7A63 <cjk>
	0x8FF6: '蒸' // U+84B8 <cjk>
	0x8FF7: '譲' // U+8B72 <cjk>
	0x8FF8: '醸' // U+91B8 <cjk>
	0x8FF9: '錠' // U+9320 <cjk>
	0x8FFA: '嘱' // U+5631 <cjk>
	0x8FFB: '埴' // U+57F4 <cjk>
	0x8FFC: '飾' // U+98FE <cjk>
	0x9040: '拭' // U+62ED <cjk>
	0x9041: '植' // U+690D <cjk>
	0x9042: '殖' // U+6B96 <cjk>
	0x9043: '燭' // U+71ED <cjk>
	0x9044: '織' // U+7E54 <cjk>
	0x9045: '職' // U+8077 <cjk>
	0x9046: '色' // U+8272 <cjk>
	0x9047: '触' // U+89E6 <cjk>
	0x9048: '食' // U+98DF <cjk>
	0x9049: '蝕' // U+8755 <cjk>
	0x904A: '辱' // U+8FB1 <cjk>
	0x904B: '尻' // U+5C3B <cjk>
	0x904C: '伸' // U+4F38 <cjk>
	0x904D: '信' // U+4FE1 <cjk>
	0x904E: '侵' // U+4FB5 <cjk>
	0x904F: '唇' // U+5507 <cjk>
	0x9050: '娠' // U+5A20 <cjk>
	0x9051: '寝' // U+5BDD <cjk>
	0x9052: '審' // U+5BE9 <cjk>
	0x9053: '心' // U+5FC3 <cjk>
	0x9054: '慎' // U+614E <cjk>
	0x9055: '振' // U+632F <cjk>
	0x9056: '新' // U+65B0 <cjk>
	0x9057: '晋' // U+664B <cjk>
	0x9058: '森' // U+68EE <cjk>
	0x9059: '榛' // U+699B <cjk>
	0x905A: '浸' // U+6D78 <cjk>
	0x905B: '深' // U+6DF1 <cjk>
	0x905C: '申' // U+7533 <cjk>
	0x905D: '疹' // U+75B9 <cjk>
	0x905E: '真' // U+771F <cjk>
	0x905F: '神' // U+795E <cjk>
	0x9060: '秦' // U+79E6 <cjk>
	0x9061: '紳' // U+7D33 <cjk>
	0x9062: '臣' // U+81E3 <cjk>
	0x9063: '芯' // U+82AF <cjk>
	0x9064: '薪' // U+85AA <cjk>
	0x9065: '親' // U+89AA <cjk>
	0x9066: '診' // U+8A3A <cjk>
	0x9067: '身' // U+8EAB <cjk>
	0x9068: '辛' // U+8F9B <cjk>
	0x9069: '進' // U+9032 <cjk>
	0x906A: '針' // U+91DD <cjk>
	0x906B: '震' // U+9707 <cjk>
	0x906C: '人' // U+4EBA <cjk>
	0x906D: '仁' // U+4EC1 <cjk>
	0x906E: '刃' // U+5203 <cjk>
	0x906F: '塵' // U+5875 <cjk>
	0x9070: '壬' // U+58EC <cjk>
	0x9071: '尋' // U+5C0B <cjk>
	0x9072: '甚' // U+751A <cjk>
	0x9073: '尽' // U+5C3D <cjk>
	0x9074: '腎' // U+814E <cjk>
	0x9075: '訊' // U+8A0A <cjk>
	0x9076: '迅' // U+8FC5 <cjk>
	0x9077: '陣' // U+9663 <cjk>
	0x9078: '靭' // U+976D <cjk>
	0x9079: '笥' // U+7B25 <cjk>
	0x907A: '諏' // U+8ACF <cjk>
	0x907B: '須' // U+9808 <cjk>
	0x907C: '酢' // U+9162 <cjk>
	0x907D: '図' // U+56F3 <cjk>
	0x907E: '厨' // U+53A8 <cjk>
	0x9080: '逗' // U+9017 <cjk>
	0x9081: '吹' // U+5439 <cjk>
	0x9082: '垂' // U+5782 <cjk>
	0x9083: '帥' // U+5E25 <cjk>
	0x9084: '推' // U+63A8 <cjk>
	0x9085: '水' // U+6C34 <cjk>
	0x9086: '炊' // U+708A <cjk>
	0x9087: '睡' // U+7761 <cjk>
	0x9088: '粋' // U+7C8B <cjk>
	0x9089: '翠' // U+7FE0 <cjk>
	0x908A: '衰' // U+8870 <cjk>
	0x908B: '遂' // U+9042 <cjk>
	0x908C: '酔' // U+9154 <cjk>
	0x908D: '錐' // U+9310 <cjk>
	0x908E: '錘' // U+9318 <cjk>
	0x908F: '随' // U+968F <cjk>
	0x9090: '瑞' // U+745E <cjk>
	0x9091: '髄' // U+9AC4 <cjk>
	0x9092: '崇' // U+5D07 <cjk>
	0x9093: '嵩' // U+5D69 <cjk>
	0x9094: '数' // U+6570 <cjk>
	0x9095: '枢' // U+67A2 <cjk>
	0x9096: '趨' // U+8DA8 <cjk>
	0x9097: '雛' // U+96DB <cjk>
	0x9098: '据' // U+636E <cjk>
	0x9099: '杉' // U+6749 <cjk>
	0x909A: '椙' // U+6919 <cjk>
	0x909B: '菅' // U+83C5 <cjk>
	0x909C: '頗' // U+9817 <cjk>
	0x909D: '雀' // U+96C0 <cjk>
	0x909E: '裾' // U+88FE <cjk>
	0x909F: '澄' // U+6F84 <cjk>
	0x90A0: '摺' // U+647A <cjk>
	0x90A1: '寸' // U+5BF8 <cjk>
	0x90A2: '世' // U+4E16 <cjk>
	0x90A3: '瀬' // U+702C <cjk>
	0x90A4: '畝' // U+755D <cjk>
	0x90A5: '是' // U+662F <cjk>
	0x90A6: '凄' // U+51C4 <cjk>
	0x90A7: '制' // U+5236 <cjk>
	0x90A8: '勢' // U+52E2 <cjk>
	0x90A9: '姓' // U+59D3 <cjk>
	0x90AA: '征' // U+5F81 <cjk>
	0x90AB: '性' // U+6027 <cjk>
	0x90AC: '成' // U+6210 <cjk>
	0x90AD: '政' // U+653F <cjk>
	0x90AE: '整' // U+6574 <cjk>
	0x90AF: '星' // U+661F <cjk>
	0x90B0: '晴' // U+6674 <cjk>
	0x90B1: '棲' // U+68F2 <cjk>
	0x90B2: '栖' // U+6816 <cjk>
	0x90B3: '正' // U+6B63 <cjk>
	0x90B4: '清' // U+6E05 <cjk>
	0x90B5: '牲' // U+7272 <cjk>
	0x90B6: '生' // U+751F <cjk>
	0x90B7: '盛' // U+76DB <cjk>
	0x90B8: '精' // U+7CBE <cjk>
	0x90B9: '聖' // U+8056 <cjk>
	0x90BA: '声' // U+58F0 <cjk>
	0x90BB: '製' // U+88FD <cjk>
	0x90BC: '西' // U+897F <cjk>
	0x90BD: '誠' // U+8AA0 <cjk>
	0x90BE: '誓' // U+8A93 <cjk>
	0x90BF: '請' // U+8ACB <cjk>
	0x90C0: '逝' // U+901D <cjk>
	0x90C1: '醒' // U+9192 <cjk>
	0x90C2: '青' // U+9752 <cjk>
	0x90C3: '静' // U+9759 <cjk>
	0x90C4: '斉' // U+6589 <cjk>
	0x90C5: '税' // U+7A0E <cjk>
	0x90C6: '脆' // U+8106 <cjk>
	0x90C7: '隻' // U+96BB <cjk>
	0x90C8: '席' // U+5E2D <cjk>
	0x90C9: '惜' // U+60DC <cjk>
	0x90CA: '戚' // U+621A <cjk>
	0x90CB: '斥' // U+65A5 <cjk>
	0x90CC: '昔' // U+6614 <cjk>
	0x90CD: '析' // U+6790 <cjk>
	0x90CE: '石' // U+77F3 <cjk>
	0x90CF: '積' // U+7A4D <cjk>
	0x90D0: '籍' // U+7C4D <cjk>
	0x90D1: '績' // U+7E3E <cjk>
	0x90D2: '脊' // U+810A <cjk>
	0x90D3: '責' // U+8CAC <cjk>
	0x90D4: '赤' // U+8D64 <cjk>
	0x90D5: '跡' // U+8DE1 <cjk>
	0x90D6: '蹟' // U+8E5F <cjk>
	0x90D7: '碩' // U+78A9 <cjk>
	0x90D8: '切' // U+5207 <cjk>
	0x90D9: '拙' // U+62D9 <cjk>
	0x90DA: '接' // U+63A5 <cjk>
	0x90DB: '摂' // U+6442 <cjk>
	0x90DC: '折' // U+6298 <cjk>
	0x90DD: '設' // U+8A2D <cjk>
	0x90DE: '窃' // U+7A83 <cjk>
	0x90DF: '節' // U+7BC0 <cjk>
	0x90E0: '説' // U+8AAC <cjk>
	0x90E1: '雪' // U+96EA <cjk>
	0x90E2: '絶' // U+7D76 <cjk>
	0x90E3: '舌' // U+820C <cjk>
	0x90E4: '蝉' // U+8749 <cjk>
	0x90E5: '仙' // U+4ED9 <cjk>
	0x90E6: '先' // U+5148 <cjk>
	0x90E7: '千' // U+5343 <cjk>
	0x90E8: '占' // U+5360 <cjk>
	0x90E9: '宣' // U+5BA3 <cjk>
	0x90EA: '専' // U+5C02 <cjk>
	0x90EB: '尖' // U+5C16 <cjk>
	0x90EC: '川' // U+5DDD <cjk>
	0x90ED: '戦' // U+6226 <cjk>
	0x90EE: '扇' // U+6247 <cjk>
	0x90EF: '撰' // U+64B0 <cjk>
	0x90F0: '栓' // U+6813 <cjk>
	0x90F1: '栴' // U+6834 <cjk>
	0x90F2: '泉' // U+6CC9 <cjk>
	0x90F3: '浅' // U+6D45 <cjk>
	0x90F4: '洗' // U+6D17 <cjk>
	0x90F5: '染' // U+67D3 <cjk>
	0x90F6: '潜' // U+6F5C <cjk>
	0x90F7: '煎' // U+714E <cjk>
	0x90F8: '煽' // U+717D <cjk>
	0x90F9: '旋' // U+65CB <cjk>
	0x90FA: '穿' // U+7A7F <cjk>
	0x90FB: '箭' // U+7BAD <cjk>
	0x90FC: '線' // U+7DDA <cjk>
	0x9140: '繊' // U+7E4A <cjk>
	0x9141: '羨' // U+7FA8 <cjk>
	0x9142: '腺' // U+817A <cjk>
	0x9143: '舛' // U+821B <cjk>
	0x9144: '船' // U+8239 <cjk>
	0x9145: '薦' // U+85A6 <cjk>
	0x9146: '詮' // U+8A6E <cjk>
	0x9147: '賎' // U+8CCE <cjk>
	0x9148: '践' // U+8DF5 <cjk>
	0x9149: '選' // U+9078 <cjk>
	0x914A: '遷' // U+9077 <cjk>
	0x914B: '銭' // U+92AD <cjk>
	0x914C: '銑' // U+9291 <cjk>
	0x914D: '閃' // U+9583 <cjk>
	0x914E: '鮮' // U+9BAE <cjk>
	0x914F: '前' // U+524D <cjk>
	0x9150: '善' // U+5584 <cjk>
	0x9151: '漸' // U+6F38 <cjk>
	0x9152: '然' // U+7136 <cjk>
	0x9153: '全' // U+5168 <cjk>
	0x9154: '禅' // U+7985 <cjk>
	0x9155: '繕' // U+7E55 <cjk>
	0x9156: '膳' // U+81B3 <cjk>
	0x9157: '糎' // U+7CCE <cjk>
	0x9158: '噌' // U+564C <cjk>
	0x9159: '塑' // U+5851 <cjk>
	0x915A: '岨' // U+5CA8 <cjk>
	0x915B: '措' // U+63AA <cjk>
	0x915C: '曾' // U+66FE <cjk>
	0x915D: '曽' // U+66FD <cjk>
	0x915E: '楚' // U+695A <cjk>
	0x915F: '狙' // U+72D9 <cjk>
	0x9160: '疏' // U+758F <cjk>
	0x9161: '疎' // U+758E <cjk>
	0x9162: '礎' // U+790E <cjk>
	0x9163: '祖' // U+7956 <cjk>
	0x9164: '租' // U+79DF <cjk>
	0x9165: '粗' // U+7C97 <cjk>
	0x9166: '素' // U+7D20 <cjk>
	0x9167: '組' // U+7D44 <cjk>
	0x9168: '蘇' // U+8607 <cjk>
	0x9169: '訴' // U+8A34 <cjk>
	0x916A: '阻' // U+963B <cjk>
	0x916B: '遡' // U+9061 <cjk>
	0x916C: '鼠' // U+9F20 <cjk>
	0x916D: '僧' // U+50E7 <cjk>
	0x916E: '創' // U+5275 <cjk>
	0x916F: '双' // U+53CC <cjk>
	0x9170: '叢' // U+53E2 <cjk>
	0x9171: '倉' // U+5009 <cjk>
	0x9172: '喪' // U+55AA <cjk>
	0x9173: '壮' // U+58EE <cjk>
	0x9174: '奏' // U+594F <cjk>
	0x9175: '爽' // U+723D <cjk>
	0x9176: '宋' // U+5B8B <cjk>
	0x9177: '層' // U+5C64 <cjk>
	0x9178: '匝' // U+531D <cjk>
	0x9179: '惣' // U+60E3 <cjk>
	0x917A: '想' // U+60F3 <cjk>
	0x917B: '捜' // U+635C <cjk>
	0x917C: '掃' // U+6383 <cjk>
	0x917D: '挿' // U+633F <cjk>
	0x917E: '掻' // U+63BB <cjk>
	0x9180: '操' // U+64CD <cjk>
	0x9181: '早' // U+65E9 <cjk>
	0x9182: '曹' // U+66F9 <cjk>
	0x9183: '巣' // U+5DE3 <cjk>
	0x9184: '槍' // U+69CD <cjk>
	0x9185: '槽' // U+69FD <cjk>
	0x9186: '漕' // U+6F15 <cjk>
	0x9187: '燥' // U+71E5 <cjk>
	0x9188: '争' // U+4E89 <cjk>
	0x9189: '痩' // U+75E9 <cjk>
	0x918A: '相' // U+76F8 <cjk>
	0x918B: '窓' // U+7A93 <cjk>
	0x918C: '糟' // U+7CDF <cjk>
	0x918D: '総' // U+7DCF <cjk>
	0x918E: '綜' // U+7D9C <cjk>
	0x918F: '聡' // U+8061 <cjk>
	0x9190: '草' // U+8349 <cjk>
	0x9191: '荘' // U+8358 <cjk>
	0x9192: '葬' // U+846C <cjk>
	0x9193: '蒼' // U+84BC <cjk>
	0x9194: '藻' // U+85FB <cjk>
	0x9195: '装' // U+88C5 <cjk>
	0x9196: '走' // U+8D70 <cjk>
	0x9197: '送' // U+9001 <cjk>
	0x9198: '遭' // U+906D <cjk>
	0x9199: '鎗' // U+9397 <cjk>
	0x919A: '霜' // U+971C <cjk>
	0x919B: '騒' // U+9A12 <cjk>
	0x919C: '像' // U+50CF <cjk>
	0x919D: '増' // U+5897 <cjk>
	0x919E: '憎' // U+618E <cjk>
	0x919F: '臓' // U+81D3 <cjk>
	0x91A0: '蔵' // U+8535 <cjk>
	0x91A1: '贈' // U+8D08 <cjk>
	0x91A2: '造' // U+9020 <cjk>
	0x91A3: '促' // U+4FC3 <cjk>
	0x91A4: '側' // U+5074 <cjk>
	0x91A5: '則' // U+5247 <cjk>
	0x91A6: '即' // U+5373 <cjk>
	0x91A7: '息' // U+606F <cjk>
	0x91A8: '捉' // U+6349 <cjk>
	0x91A9: '束' // U+675F <cjk>
	0x91AA: '測' // U+6E2C <cjk>
	0x91AB: '足' // U+8DB3 <cjk>
	0x91AC: '速' // U+901F <cjk>
	0x91AD: '俗' // U+4FD7 <cjk>
	0x91AE: '属' // U+5C5E <cjk>
	0x91AF: '賊' // U+8CCA <cjk>
	0x91B0: '族' // U+65CF <cjk>
	0x91B1: '続' // U+7D9A <cjk>
	0x91B2: '卒' // U+5352 <cjk>
	0x91B3: '袖' // U+8896 <cjk>
	0x91B4: '其' // U+5176 <cjk>
	0x91B5: '揃' // U+63C3 <cjk>
	0x91B6: '存' // U+5B58 <cjk>
	0x91B7: '孫' // U+5B6B <cjk>
	0x91B8: '尊' // U+5C0A <cjk>
	0x91B9: '損' // U+640D <cjk>
	0x91BA: '村' // U+6751 <cjk>
	0x91BB: '遜' // U+905C <cjk>
	0x91BC: '他' // U+4ED6 <cjk>
	0x91BD: '多' // U+591A <cjk>
	0x91BE: '太' // U+592A <cjk>
	0x91BF: '汰' // U+6C70 <cjk>
	0x91C0: '詑' // U+8A51 <cjk>
	0x91C1: '唾' // U+553E <cjk>
	0x91C2: '堕' // U+5815 <cjk>
	0x91C3: '妥' // U+59A5 <cjk>
	0x91C4: '惰' // U+60F0 <cjk>
	0x91C5: '打' // U+6253 <cjk>
	0x91C6: '柁' // U+67C1 <cjk>
	0x91C7: '舵' // U+8235 <cjk>
	0x91C8: '楕' // U+6955 <cjk>
	0x91C9: '陀' // U+9640 <cjk>
	0x91CA: '駄' // U+99C4 <cjk>
	0x91CB: '騨' // U+9A28 <cjk>
	0x91CC: '体' // U+4F53 <cjk>
	0x91CD: '堆' // U+5806 <cjk>
	0x91CE: '対' // U+5BFE <cjk>
	0x91CF: '耐' // U+8010 <cjk>
	0x91D0: '岱' // U+5CB1 <cjk>
	0x91D1: '帯' // U+5E2F <cjk>
	0x91D2: '待' // U+5F85 <cjk>
	0x91D3: '怠' // U+6020 <cjk>
	0x91D4: '態' // U+614B <cjk>
	0x91D5: '戴' // U+6234 <cjk>
	0x91D6: '替' // U+66FF <cjk>
	0x91D7: '泰' // U+6CF0 <cjk>
	0x91D8: '滞' // U+6EDE <cjk>
	0x91D9: '胎' // U+80CE <cjk>
	0x91DA: '腿' // U+817F <cjk>
	0x91DB: '苔' // U+82D4 <cjk>
	0x91DC: '袋' // U+888B <cjk>
	0x91DD: '貸' // U+8CB8 <cjk>
	0x91DE: '退' // U+9000 <cjk>
	0x91DF: '逮' // U+902E <cjk>
	0x91E0: '隊' // U+968A <cjk>
	0x91E1: '黛' // U+9EDB <cjk>
	0x91E2: '鯛' // U+9BDB <cjk>
	0x91E3: '代' // U+4EE3 <cjk>
	0x91E4: '台' // U+53F0 <cjk>
	0x91E5: '大' // U+5927 <cjk>
	0x91E6: '第' // U+7B2C <cjk>
	0x91E7: '醍' // U+918D <cjk>
	0x91E8: '題' // U+984C <cjk>
	0x91E9: '鷹' // U+9DF9 <cjk>
	0x91EA: '滝' // U+6EDD <cjk>
	0x91EB: '瀧' // U+7027 <cjk>
	0x91EC: '卓' // U+5353 <cjk>
	0x91ED: '啄' // U+5544 <cjk>
	0x91EE: '宅' // U+5B85 <cjk>
	0x91EF: '托' // U+6258 <cjk>
	0x91F0: '択' // U+629E <cjk>
	0x91F1: '拓' // U+62D3 <cjk>
	0x91F2: '沢' // U+6CA2 <cjk>
	0x91F3: '濯' // U+6FEF <cjk>
	0x91F4: '琢' // U+7422 <cjk>
	0x91F5: '託' // U+8A17 <cjk>
	0x91F6: '鐸' // U+9438 <cjk>
	0x91F7: '濁' // U+6FC1 <cjk>
	0x91F8: '諾' // U+8AFE <cjk>
	0x91F9: '茸' // U+8338 <cjk>
	0x91FA: '凧' // U+51E7 <cjk>
	0x91FB: '蛸' // U+86F8 <cjk>
	0x91FC: '只' // U+53EA <cjk>
	0x9240: '叩' // U+53E9 <cjk>
	0x9241: '但' // U+4F46 <cjk>
	0x9242: '達' // U+9054 <cjk>
	0x9243: '辰' // U+8FB0 <cjk>
	0x9244: '奪' // U+596A <cjk>
	0x9245: '脱' // U+8131 <cjk>
	0x9246: '巽' // U+5DFD <cjk>
	0x9247: '竪' // U+7AEA <cjk>
	0x9248: '辿' // U+8FBF <cjk>
	0x9249: '棚' // U+68DA <cjk>
	0x924A: '谷' // U+8C37 <cjk>
	0x924B: '狸' // U+72F8 <cjk>
	0x924C: '鱈' // U+9C48 <cjk>
	0x924D: '樽' // U+6A3D <cjk>
	0x924E: '誰' // U+8AB0 <cjk>
	0x924F: '丹' // U+4E39 <cjk>
	0x9250: '単' // U+5358 <cjk>
	0x9251: '嘆' // U+5606 <cjk>
	0x9252: '坦' // U+5766 <cjk>
	0x9253: '担' // U+62C5 <cjk>
	0x9254: '探' // U+63A2 <cjk>
	0x9255: '旦' // U+65E6 <cjk>
	0x9256: '歎' // U+6B4E <cjk>
	0x9257: '淡' // U+6DE1 <cjk>
	0x9258: '湛' // U+6E5B <cjk>
	0x9259: '炭' // U+70AD <cjk>
	0x925A: '短' // U+77ED <cjk>
	0x925B: '端' // U+7AEF <cjk>
	0x925C: '箪' // U+7BAA <cjk>
	0x925D: '綻' // U+7DBB <cjk>
	0x925E: '耽' // U+803D <cjk>
	0x925F: '胆' // U+80C6 <cjk>
	0x9260: '蛋' // U+86CB <cjk>
	0x9261: '誕' // U+8A95 <cjk>
	0x9262: '鍛' // U+935B <cjk>
	0x9263: '団' // U+56E3 <cjk>
	0x9264: '壇' // U+58C7 <cjk>
	0x9265: '弾' // U+5F3E <cjk>
	0x9266: '断' // U+65AD <cjk>
	0x9267: '暖' // U+6696 <cjk>
	0x9268: '檀' // U+6A80 <cjk>
	0x9269: '段' // U+6BB5 <cjk>
	0x926A: '男' // U+7537 <cjk>
	0x926B: '談' // U+8AC7 <cjk>
	0x926C: '値' // U+5024 <cjk>
	0x926D: '知' // U+77E5 <cjk>
	0x926E: '地' // U+5730 <cjk>
	0x926F: '弛' // U+5F1B <cjk>
	0x9270: '恥' // U+6065 <cjk>
	0x9271: '智' // U+667A <cjk>
	0x9272: '池' // U+6C60 <cjk>
	0x9273: '痴' // U+75F4 <cjk>
	0x9274: '稚' // U+7A1A <cjk>
	0x9275: '置' // U+7F6E <cjk>
	0x9276: '致' // U+81F4 <cjk>
	0x9277: '蜘' // U+8718 <cjk>
	0x9278: '遅' // U+9045 <cjk>
	0x9279: '馳' // U+99B3 <cjk>
	0x927A: '築' // U+7BC9 <cjk>
	0x927B: '畜' // U+755C <cjk>
	0x927C: '竹' // U+7AF9 <cjk>
	0x927D: '筑' // U+7B51 <cjk>
	0x927E: '蓄' // U+84C4 <cjk>
	0x9280: '逐' // U+9010 <cjk>
	0x9281: '秩' // U+79E9 <cjk>
	0x9282: '窒' // U+7A92 <cjk>
	0x9283: '茶' // U+8336 <cjk>
	0x9284: '嫡' // U+5AE1 <cjk>
	0x9285: '着' // U+7740 <cjk>
	0x9286: '中' // U+4E2D <cjk>
	0x9287: '仲' // U+4EF2 <cjk>
	0x9288: '宙' // U+5B99 <cjk>
	0x9289: '忠' // U+5FE0 <cjk>
	0x928A: '抽' // U+62BD <cjk>
	0x928B: '昼' // U+663C <cjk>
	0x928C: '柱' // U+67F1 <cjk>
	0x928D: '注' // U+6CE8 <cjk>
	0x928E: '虫' // U+866B <cjk>
	0x928F: '衷' // U+8877 <cjk>
	0x9290: '註' // U+8A3B <cjk>
	0x9291: '酎' // U+914E <cjk>
	0x9292: '鋳' // U+92F3 <cjk>
	0x9293: '駐' // U+99D0 <cjk>
	0x9294: '樗' // U+6A17 <cjk>
	0x9295: '瀦' // U+7026 <cjk>
	0x9296: '猪' // U+732A <cjk>
	0x9297: '苧' // U+82E7 <cjk>
	0x9298: '著' // U+8457 <cjk>
	0x9299: '貯' // U+8CAF <cjk>
	0x929A: '丁' // U+4E01 <cjk>
	0x929B: '兆' // U+5146 <cjk>
	0x929C: '凋' // U+51CB <cjk>
	0x929D: '喋' // U+558B <cjk>
	0x929E: '寵' // U+5BF5 <cjk>
	0x929F: '帖' // U+5E16 <cjk>
	0x92A0: '帳' // U+5E33 <cjk>
	0x92A1: '庁' // U+5E81 <cjk>
	0x92A2: '弔' // U+5F14 <cjk>
	0x92A3: '張' // U+5F35 <cjk>
	0x92A4: '彫' // U+5F6B <cjk>
	0x92A5: '徴' // U+5FB4 <cjk>
	0x92A6: '懲' // U+61F2 <cjk>
	0x92A7: '挑' // U+6311 <cjk>
	0x92A8: '暢' // U+66A2 <cjk>
	0x92A9: '朝' // U+671D <cjk>
	0x92AA: '潮' // U+6F6E <cjk>
	0x92AB: '牒' // U+7252 <cjk>
	0x92AC: '町' // U+753A <cjk>
	0x92AD: '眺' // U+773A <cjk>
	0x92AE: '聴' // U+8074 <cjk>
	0x92AF: '脹' // U+8139 <cjk>
	0x92B0: '腸' // U+8178 <cjk>
	0x92B1: '蝶' // U+8776 <cjk>
	0x92B2: '調' // U+8ABF <cjk>
	0x92B3: '諜' // U+8ADC <cjk>
	0x92B4: '超' // U+8D85 <cjk>
	0x92B5: '跳' // U+8DF3 <cjk>
	0x92B6: '銚' // U+929A <cjk>
	0x92B7: '長' // U+9577 <cjk>
	0x92B8: '頂' // U+9802 <cjk>
	0x92B9: '鳥' // U+9CE5 <cjk>
	0x92BA: '勅' // U+52C5 <cjk>
	0x92BB: '捗' // U+6357 <cjk>
	0x92BC: '直' // U+76F4 <cjk>
	0x92BD: '朕' // U+6715 <cjk>
	0x92BE: '沈' // U+6C88 <cjk>
	0x92BF: '珍' // U+73CD <cjk>
	0x92C0: '賃' // U+8CC3 <cjk>
	0x92C1: '鎮' // U+93AE <cjk>
	0x92C2: '陳' // U+9673 <cjk>
	0x92C3: '津' // U+6D25 <cjk>
	0x92C4: '墜' // U+589C <cjk>
	0x92C5: '椎' // U+690E <cjk>
	0x92C6: '槌' // U+69CC <cjk>
	0x92C7: '追' // U+8FFD <cjk>
	0x92C8: '鎚' // U+939A <cjk>
	0x92C9: '痛' // U+75DB <cjk>
	0x92CA: '通' // U+901A <cjk>
	0x92CB: '塚' // U+585A <cjk>
	0x92CC: '栂' // U+6802 <cjk>
	0x92CD: '掴' // U+63B4 <cjk>
	0x92CE: '槻' // U+69FB <cjk>
	0x92CF: '佃' // U+4F43 <cjk>
	0x92D0: '漬' // U+6F2C <cjk>
	0x92D1: '柘' // U+67D8 <cjk>
	0x92D2: '辻' // U+8FBB <cjk>
	0x92D3: '蔦' // U+8526 <cjk>
	0x92D4: '綴' // U+7DB4 <cjk>
	0x92D5: '鍔' // U+9354 <cjk>
	0x92D6: '椿' // U+693F <cjk>
	0x92D7: '潰' // U+6F70 <cjk>
	0x92D8: '坪' // U+576A <cjk>
	0x92D9: '壷' // U+58F7 <cjk>
	0x92DA: '嬬' // U+5B2C <cjk>
	0x92DB: '紬' // U+7D2C <cjk>
	0x92DC: '爪' // U+722A <cjk>
	0x92DD: '吊' // U+540A <cjk>
	0x92DE: '釣' // U+91E3 <cjk>
	0x92DF: '鶴' // U+9DB4 <cjk>
	0x92E0: '亭' // U+4EAD <cjk>
	0x92E1: '低' // U+4F4E <cjk>
	0x92E2: '停' // U+505C <cjk>
	0x92E3: '偵' // U+5075 <cjk>
	0x92E4: '剃' // U+5243 <cjk>
	0x92E5: '貞' // U+8C9E <cjk>
	0x92E6: '呈' // U+5448 <cjk>
	0x92E7: '堤' // U+5824 <cjk>
	0x92E8: '定' // U+5B9A <cjk>
	0x92E9: '帝' // U+5E1D <cjk>
	0x92EA: '底' // U+5E95 <cjk>
	0x92EB: '庭' // U+5EAD <cjk>
	0x92EC: '廷' // U+5EF7 <cjk>
	0x92ED: '弟' // U+5F1F <cjk>
	0x92EE: '悌' // U+608C <cjk>
	0x92EF: '抵' // U+62B5 <cjk>
	0x92F0: '挺' // U+633A <cjk>
	0x92F1: '提' // U+63D0 <cjk>
	0x92F2: '梯' // U+68AF <cjk>
	0x92F3: '汀' // U+6C40 <cjk>
	0x92F4: '碇' // U+7887 <cjk>
	0x92F5: '禎' // U+798E <cjk>
	0x92F6: '程' // U+7A0B <cjk>
	0x92F7: '締' // U+7DE0 <cjk>
	0x92F8: '艇' // U+8247 <cjk>
	0x92F9: '訂' // U+8A02 <cjk>
	0x92FA: '諦' // U+8AE6 <cjk>
	0x92FB: '蹄' // U+8E44 <cjk>
	0x92FC: '逓' // U+9013 <cjk>
	0x9340: '邸' // U+90B8 <cjk>
	0x9341: '鄭' // U+912D <cjk>
	0x9342: '釘' // U+91D8 <cjk>
	0x9343: '鼎' // U+9F0E <cjk>
	0x9344: '泥' // U+6CE5 <cjk>
	0x9345: '摘' // U+6458 <cjk>
	0x9346: '擢' // U+64E2 <cjk>
	0x9347: '敵' // U+6575 <cjk>
	0x9348: '滴' // U+6EF4 <cjk>
	0x9349: '的' // U+7684 <cjk>
	0x934A: '笛' // U+7B1B <cjk>
	0x934B: '適' // U+9069 <cjk>
	0x934C: '鏑' // U+93D1 <cjk>
	0x934D: '溺' // U+6EBA <cjk>
	0x934E: '哲' // U+54F2 <cjk>
	0x934F: '徹' // U+5FB9 <cjk>
	0x9350: '撤' // U+64A4 <cjk>
	0x9351: '轍' // U+8F4D <cjk>
	0x9352: '迭' // U+8FED <cjk>
	0x9353: '鉄' // U+9244 <cjk>
	0x9354: '典' // U+5178 <cjk>
	0x9355: '填' // U+586B <cjk>
	0x9356: '天' // U+5929 <cjk>
	0x9357: '展' // U+5C55 <cjk>
	0x9358: '店' // U+5E97 <cjk>
	0x9359: '添' // U+6DFB <cjk>
	0x935A: '纏' // U+7E8F <cjk>
	0x935B: '甜' // U+751C <cjk>
	0x935C: '貼' // U+8CBC <cjk>
	0x935D: '転' // U+8EE2 <cjk>
	0x935E: '顛' // U+985B <cjk>
	0x935F: '点' // U+70B9 <cjk>
	0x9360: '伝' // U+4F1D <cjk>
	0x9361: '殿' // U+6BBF <cjk>
	0x9362: '澱' // U+6FB1 <cjk>
	0x9363: '田' // U+7530 <cjk>
	0x9364: '電' // U+96FB <cjk>
	0x9365: '兎' // U+514E <cjk>
	0x9366: '吐' // U+5410 <cjk>
	0x9367: '堵' // U+5835 <cjk>
	0x9368: '塗' // U+5857 <cjk>
	0x9369: '妬' // U+59AC <cjk>
	0x936A: '屠' // U+5C60 <cjk>
	0x936B: '徒' // U+5F92 <cjk>
	0x936C: '斗' // U+6597 <cjk>
	0x936D: '杜' // U+675C <cjk>
	0x936E: '渡' // U+6E21 <cjk>
	0x936F: '登' // U+767B <cjk>
	0x9370: '菟' // U+83DF <cjk>
	0x9371: '賭' // U+8CED <cjk>
	0x9372: '途' // U+9014 <cjk>
	0x9373: '都' // U+90FD <cjk>
	0x9374: '鍍' // U+934D <cjk>
	0x9375: '砥' // U+7825 <cjk>
	0x9376: '砺' // U+783A <cjk>
	0x9377: '努' // U+52AA <cjk>
	0x9378: '度' // U+5EA6 <cjk>
	0x9379: '土' // U+571F <cjk>
	0x937A: '奴' // U+5974 <cjk>
	0x937B: '怒' // U+6012 <cjk>
	0x937C: '倒' // U+5012 <cjk>
	0x937D: '党' // U+515A <cjk>
	0x937E: '冬' // U+51AC <cjk>
	0x9380: '凍' // U+51CD <cjk>
	0x9381: '刀' // U+5200 <cjk>
	0x9382: '唐' // U+5510 <cjk>
	0x9383: '塔' // U+5854 <cjk>
	0x9384: '塘' // U+5858 <cjk>
	0x9385: '套' // U+5957 <cjk>
	0x9386: '宕' // U+5B95 <cjk>
	0x9387: '島' // U+5CF6 <cjk>
	0x9388: '嶋' // U+5D8B <cjk>
	0x9389: '悼' // U+60BC <cjk>
	0x938A: '投' // U+6295 <cjk>
	0x938B: '搭' // U+642D <cjk>
	0x938C: '東' // U+6771 <cjk>
	0x938D: '桃' // U+6843 <cjk>
	0x938E: '梼' // U+68BC <cjk>
	0x938F: '棟' // U+68DF <cjk>
	0x9390: '盗' // U+76D7 <cjk>
	0x9391: '淘' // U+6DD8 <cjk>
	0x9392: '湯' // U+6E6F <cjk>
	0x9393: '涛' // U+6D9B <cjk>
	0x9394: '灯' // U+706F <cjk>
	0x9395: '燈' // U+71C8 <cjk>
	0x9396: '当' // U+5F53 <cjk>
	0x9397: '痘' // U+75D8 <cjk>
	0x9398: '祷' // U+7977 <cjk>
	0x9399: '等' // U+7B49 <cjk>
	0x939A: '答' // U+7B54 <cjk>
	0x939B: '筒' // U+7B52 <cjk>
	0x939C: '糖' // U+7CD6 <cjk>
	0x939D: '統' // U+7D71 <cjk>
	0x939E: '到' // U+5230 <cjk>
	0x939F: '董' // U+8463 <cjk>
	0x93A0: '蕩' // U+8569 <cjk>
	0x93A1: '藤' // U+85E4 <cjk>
	0x93A2: '討' // U+8A0E <cjk>
	0x93A3: '謄' // U+8B04 <cjk>
	0x93A4: '豆' // U+8C46 <cjk>
	0x93A5: '踏' // U+8E0F <cjk>
	0x93A6: '逃' // U+9003 <cjk>
	0x93A7: '透' // U+900F <cjk>
	0x93A8: '鐙' // U+9419 <cjk>
	0x93A9: '陶' // U+9676 <cjk>
	0x93AA: '頭' // U+982D <cjk>
	0x93AB: '騰' // U+9A30 <cjk>
	0x93AC: '闘' // U+95D8 <cjk>
	0x93AD: '働' // U+50CD <cjk>
	0x93AE: '動' // U+52D5 <cjk>
	0x93AF: '同' // U+540C <cjk>
	0x93B0: '堂' // U+5802 <cjk>
	0x93B1: '導' // U+5C0E <cjk>
	0x93B2: '憧' // U+61A7 <cjk>
	0x93B3: '撞' // U+649E <cjk>
	0x93B4: '洞' // U+6D1E <cjk>
	0x93B5: '瞳' // U+77B3 <cjk>
	0x93B6: '童' // U+7AE5 <cjk>
	0x93B7: '胴' // U+80F4 <cjk>
	0x93B8: '萄' // U+8404 <cjk>
	0x93B9: '道' // U+9053 <cjk>
	0x93BA: '銅' // U+9285 <cjk>
	0x93BB: '峠' // U+5CE0 <cjk>
	0x93BC: '鴇' // U+9D07 <cjk>
	0x93BD: '匿' // U+533F <cjk>
	0x93BE: '得' // U+5F97 <cjk>
	0x93BF: '徳' // U+5FB3 <cjk>
	0x93C0: '涜' // U+6D9C <cjk>
	0x93C1: '特' // U+7279 <cjk>
	0x93C2: '督' // U+7763 <cjk>
	0x93C3: '禿' // U+79BF <cjk>
	0x93C4: '篤' // U+7BE4 <cjk>
	0x93C5: '毒' // U+6BD2 <cjk>
	0x93C6: '独' // U+72EC <cjk>
	0x93C7: '読' // U+8AAD <cjk>
	0x93C8: '栃' // U+6803 <cjk>
	0x93C9: '橡' // U+6A61 <cjk>
	0x93CA: '凸' // U+51F8 <cjk>
	0x93CB: '突' // U+7A81 <cjk>
	0x93CC: '椴' // U+6934 <cjk>
	0x93CD: '届' // U+5C4A <cjk>
	0x93CE: '鳶' // U+9CF6 <cjk>
	0x93CF: '苫' // U+82EB <cjk>
	0x93D0: '寅' // U+5BC5 <cjk>
	0x93D1: '酉' // U+9149 <cjk>
	0x93D2: '瀞' // U+701E <cjk>
	0x93D3: '噸' // U+5678 <cjk>
	0x93D4: '屯' // U+5C6F <cjk>
	0x93D5: '惇' // U+60C7 <cjk>
	0x93D6: '敦' // U+6566 <cjk>
	0x93D7: '沌' // U+6C8C <cjk>
	0x93D8: '豚' // U+8C5A <cjk>
	0x93D9: '遁' // U+9041 <cjk>
	0x93DA: '頓' // U+9813 <cjk>
	0x93DB: '呑' // U+5451 <cjk>
	0x93DC: '曇' // U+66C7 <cjk>
	0x93DD: '鈍' // U+920D <cjk>
	0x93DE: '奈' // U+5948 <cjk>
	0x93DF: '那' // U+90A3 <cjk>
	0x93E0: '内' // U+5185 <cjk>
	0x93E1: '乍' // U+4E4D <cjk>
	0x93E2: '凪' // U+51EA <cjk>
	0x93E3: '薙' // U+8599 <cjk>
	0x93E4: '謎' // U+8B0E <cjk>
	0x93E5: '灘' // U+7058 <cjk>
	0x93E6: '捺' // U+637A <cjk>
	0x93E7: '鍋' // U+934B <cjk>
	0x93E8: '楢' // U+6962 <cjk>
	0x93E9: '馴' // U+99B4 <cjk>
	0x93EA: '縄' // U+7E04 <cjk>
	0x93EB: '畷' // U+7577 <cjk>
	0x93EC: '南' // U+5357 <cjk>
	0x93ED: '楠' // U+6960 <cjk>
	0x93EE: '軟' // U+8EDF <cjk>
	0x93EF: '難' // U+96E3 <cjk>
	0x93F0: '汝' // U+6C5D <cjk>
	0x93F1: '二' // U+4E8C <cjk>
	0x93F2: '尼' // U+5C3C <cjk>
	0x93F3: '弐' // U+5F10 <cjk>
	0x93F4: '迩' // U+8FE9 <cjk>
	0x93F5: '匂' // U+5302 <cjk>
	0x93F6: '賑' // U+8CD1 <cjk>
	0x93F7: '肉' // U+8089 <cjk>
	0x93F8: '虹' // U+8679 <cjk>
	0x93F9: '廿' // U+5EFF <cjk>
	0x93FA: '日' // U+65E5 <cjk>
	0x93FB: '乳' // U+4E73 <cjk>
	0x93FC: '入' // U+5165 <cjk>
	0x9440: '如' // U+5982 <cjk>
	0x9441: '尿' // U+5C3F <cjk>
	0x9442: '韮' // U+97EE <cjk>
	0x9443: '任' // U+4EFB <cjk>
	0x9444: '妊' // U+598A <cjk>
	0x9445: '忍' // U+5FCD <cjk>
	0x9446: '認' // U+8A8D <cjk>
	0x9447: '濡' // U+6FE1 <cjk>
	0x9448: '禰' // U+79B0 <cjk>
	0x9449: '祢' // U+7962 <cjk>
	0x944A: '寧' // U+5BE7 <cjk>
	0x944B: '葱' // U+8471 <cjk>
	0x944C: '猫' // U+732B <cjk>
	0x944D: '熱' // U+71B1 <cjk>
	0x944E: '年' // U+5E74 <cjk>
	0x944F: '念' // U+5FF5 <cjk>
	0x9450: '捻' // U+637B <cjk>
	0x9451: '撚' // U+649A <cjk>
	0x9452: '燃' // U+71C3 <cjk>
	0x9453: '粘' // U+7C98 <cjk>
	0x9454: '乃' // U+4E43 <cjk>
	0x9455: '廼' // U+5EFC <cjk>
	0x9456: '之' // U+4E4B <cjk>
	0x9457: '埜' // U+57DC <cjk>
	0x9458: '嚢' // U+56A2 <cjk>
	0x9459: '悩' // U+60A9 <cjk>
	0x945A: '濃' // U+6FC3 <cjk>
	0x945B: '納' // U+7D0D <cjk>
	0x945C: '能' // U+80FD <cjk>
	0x945D: '脳' // U+8133 <cjk>
	0x945E: '膿' // U+81BF <cjk>
	0x945F: '農' // U+8FB2 <cjk>
	0x9460: '覗' // U+8997 <cjk>
	0x9461: '蚤' // U+86A4 <cjk>
	0x9462: '巴' // U+5DF4 <cjk>
	0x9463: '把' // U+628A <cjk>
	0x9464: '播' // U+64AD <cjk>
	0x9465: '覇' // U+8987 <cjk>
	0x9466: '杷' // U+6777 <cjk>
	0x9467: '波' // U+6CE2 <cjk>
	0x9468: '派' // U+6D3E <cjk>
	0x9469: '琶' // U+7436 <cjk>
	0x946A: '破' // U+7834 <cjk>
	0x946B: '婆' // U+5A46 <cjk>
	0x946C: '罵' // U+7F75 <cjk>
	0x946D: '芭' // U+82AD <cjk>
	0x946E: '馬' // U+99AC <cjk>
	0x946F: '俳' // U+4FF3 <cjk>
	0x9470: '廃' // U+5EC3 <cjk>
	0x9471: '拝' // U+62DD <cjk>
	0x9472: '排' // U+6392 <cjk>
	0x9473: '敗' // U+6557 <cjk>
	0x9474: '杯' // U+676F <cjk>
	0x9475: '盃' // U+76C3 <cjk>
	0x9476: '牌' // U+724C <cjk>
	0x9477: '背' // U+80CC <cjk>
	0x9478: '肺' // U+80BA <cjk>
	0x9479: '輩' // U+8F29 <cjk>
	0x947A: '配' // U+914D <cjk>
	0x947B: '倍' // U+500D <cjk>
	0x947C: '培' // U+57F9 <cjk>
	0x947D: '媒' // U+5A92 <cjk>
	0x947E: '梅' // U+6885 <cjk>
	0x9480: '楳' // U+6973 <cjk>
	0x9481: '煤' // U+7164 <cjk>
	0x9482: '狽' // U+72FD <cjk>
	0x9483: '買' // U+8CB7 <cjk>
	0x9484: '売' // U+58F2 <cjk>
	0x9485: '賠' // U+8CE0 <cjk>
	0x9486: '陪' // U+966A <cjk>
	0x9487: '這' // U+9019 <cjk>
	0x9488: '蝿' // U+877F <cjk>
	0x9489: '秤' // U+79E4 <cjk>
	0x948A: '矧' // U+77E7 <cjk>
	0x948B: '萩' // U+8429 <cjk>
	0x948C: '伯' // U+4F2F <cjk>
	0x948D: '剥' // U+5265 <cjk>
	0x948E: '博' // U+535A <cjk>
	0x948F: '拍' // U+62CD <cjk>
	0x9490: '柏' // U+67CF <cjk>
	0x9491: '泊' // U+6CCA <cjk>
	0x9492: '白' // U+767D <cjk>
	0x9493: '箔' // U+7B94 <cjk>
	0x9494: '粕' // U+7C95 <cjk>
	0x9495: '舶' // U+8236 <cjk>
	0x9496: '薄' // U+8584 <cjk>
	0x9497: '迫' // U+8FEB <cjk>
	0x9498: '曝' // U+66DD <cjk>
	0x9499: '漠' // U+6F20 <cjk>
	0x949A: '爆' // U+7206 <cjk>
	0x949B: '縛' // U+7E1B <cjk>
	0x949C: '莫' // U+83AB <cjk>
	0x949D: '駁' // U+99C1 <cjk>
	0x949E: '麦' // U+9EA6 <cjk>
	0x949F: '函' // U+51FD <cjk>
	0x94A0: '箱' // U+7BB1 <cjk>
	0x94A1: '硲' // U+7872 <cjk>
	0x94A2: '箸' // U+7BB8 <cjk>
	0x94A3: '肇' // U+8087 <cjk>
	0x94A4: '筈' // U+7B48 <cjk>
	0x94A5: '櫨' // U+6AE8 <cjk>
	0x94A6: '幡' // U+5E61 <cjk>
	0x94A7: '肌' // U+808C <cjk>
	0x94A8: '畑' // U+7551 <cjk>
	0x94A9: '畠' // U+7560 <cjk>
	0x94AA: '八' // U+516B <cjk>
	0x94AB: '鉢' // U+9262 <cjk>
	0x94AC: '溌' // U+6E8C <cjk>
	0x94AD: '発' // U+767A <cjk>
	0x94AE: '醗' // U+9197 <cjk>
	0x94AF: '髪' // U+9AEA <cjk>
	0x94B0: '伐' // U+4F10 <cjk>
	0x94B1: '罰' // U+7F70 <cjk>
	0x94B2: '抜' // U+629C <cjk>
	0x94B3: '筏' // U+7B4F <cjk>
	0x94B4: '閥' // U+95A5 <cjk>
	0x94B5: '鳩' // U+9CE9 <cjk>
	0x94B6: '噺' // U+567A <cjk>
	0x94B7: '塙' // U+5859 <cjk>
	0x94B8: '蛤' // U+86E4 <cjk>
	0x94B9: '隼' // U+96BC <cjk>
	0x94BA: '伴' // U+4F34 <cjk>
	0x94BB: '判' // U+5224 <cjk>
	0x94BC: '半' // U+534A <cjk>
	0x94BD: '反' // U+53CD <cjk>
	0x94BE: '叛' // U+53DB <cjk>
	0x94BF: '帆' // U+5E06 <cjk>
	0x94C0: '搬' // U+642C <cjk>
	0x94C1: '斑' // U+6591 <cjk>
	0x94C2: '板' // U+677F <cjk>
	0x94C3: '氾' // U+6C3E <cjk>
	0x94C4: '汎' // U+6C4E <cjk>
	0x94C5: '版' // U+7248 <cjk>
	0x94C6: '犯' // U+72AF <cjk>
	0x94C7: '班' // U+73ED <cjk>
	0x94C8: '畔' // U+7554 <cjk>
	0x94C9: '繁' // U+7E41 <cjk>
	0x94CA: '般' // U+822C <cjk>
	0x94CB: '藩' // U+85E9 <cjk>
	0x94CC: '販' // U+8CA9 <cjk>
	0x94CD: '範' // U+7BC4 <cjk>
	0x94CE: '釆' // U+91C6 <cjk>
	0x94CF: '煩' // U+7169 <cjk>
	0x94D0: '頒' // U+9812 <cjk>
	0x94D1: '飯' // U+98EF <cjk>
	0x94D2: '挽' // U+633D <cjk>
	0x94D3: '晩' // U+6669 <cjk>
	0x94D4: '番' // U+756A <cjk>
	0x94D5: '盤' // U+76E4 <cjk>
	0x94D6: '磐' // U+78D0 <cjk>
	0x94D7: '蕃' // U+8543 <cjk>
	0x94D8: '蛮' // U+86EE <cjk>
	0x94D9: '匪' // U+532A <cjk>
	0x94DA: '卑' // U+5351 <cjk>
	0x94DB: '否' // U+5426 <cjk>
	0x94DC: '妃' // U+5983 <cjk>
	0x94DD: '庇' // U+5E87 <cjk>
	0x94DE: '彼' // U+5F7C <cjk>
	0x94DF: '悲' // U+60B2 <cjk>
	0x94E0: '扉' // U+6249 <cjk>
	0x94E1: '批' // U+6279 <cjk>
	0x94E2: '披' // U+62AB <cjk>
	0x94E3: '斐' // U+6590 <cjk>
	0x94E4: '比' // U+6BD4 <cjk>
	0x94E5: '泌' // U+6CCC <cjk>
	0x94E6: '疲' // U+75B2 <cjk>
	0x94E7: '皮' // U+76AE <cjk>
	0x94E8: '碑' // U+7891 <cjk>
	0x94E9: '秘' // U+79D8 <cjk>
	0x94EA: '緋' // U+7DCB <cjk>
	0x94EB: '罷' // U+7F77 <cjk>
	0x94EC: '肥' // U+80A5 <cjk>
	0x94ED: '被' // U+88AB <cjk>
	0x94EE: '誹' // U+8AB9 <cjk>
	0x94EF: '費' // U+8CBB <cjk>
	0x94F0: '避' // U+907F <cjk>
	0x94F1: '非' // U+975E <cjk>
	0x94F2: '飛' // U+98DB <cjk>
	0x94F3: '樋' // U+6A0B <cjk>
	0x94F4: '簸' // U+7C38 <cjk>
	0x94F5: '備' // U+5099 <cjk>
	0x94F6: '尾' // U+5C3E <cjk>
	0x94F7: '微' // U+5FAE <cjk>
	0x94F8: '枇' // U+6787 <cjk>
	0x94F9: '毘' // U+6BD8 <cjk>
	0x94FA: '琵' // U+7435 <cjk>
	0x94FB: '眉' // U+7709 <cjk>
	0x94FC: '美' // U+7F8E <cjk>
	0x9540: '鼻' // U+9F3B <cjk>
	0x9541: '柊' // U+67CA <cjk>
	0x9542: '稗' // U+7A17 <cjk>
	0x9543: '匹' // U+5339 <cjk>
	0x9544: '疋' // U+758B <cjk>
	0x9545: '髭' // U+9AED <cjk>
	0x9546: '彦' // U+5F66 <cjk>
	0x9547: '膝' // U+819D <cjk>
	0x9548: '菱' // U+83F1 <cjk>
	0x9549: '肘' // U+8098 <cjk>
	0x954A: '弼' // U+5F3C <cjk>
	0x954B: '必' // U+5FC5 <cjk>
	0x954C: '畢' // U+7562 <cjk>
	0x954D: '筆' // U+7B46 <cjk>
	0x954E: '逼' // U+903C <cjk>
	0x954F: '桧' // U+6867 <cjk>
	0x9550: '姫' // U+59EB <cjk>
	0x9551: '媛' // U+5A9B <cjk>
	0x9552: '紐' // U+7D10 <cjk>
	0x9553: '百' // U+767E <cjk>
	0x9554: '謬' // U+8B2C <cjk>
	0x9555: '俵' // U+4FF5 <cjk>
	0x9556: '彪' // U+5F6A <cjk>
	0x9557: '標' // U+6A19 <cjk>
	0x9558: '氷' // U+6C37 <cjk>
	0x9559: '漂' // U+6F02 <cjk>
	0x955A: '瓢' // U+74E2 <cjk>
	0x955B: '票' // U+7968 <cjk>
	0x955C: '表' // U+8868 <cjk>
	0x955D: '評' // U+8A55 <cjk>
	0x955E: '豹' // U+8C79 <cjk>
	0x955F: '廟' // U+5EDF <cjk>
	0x9560: '描' // U+63CF <cjk>
	0x9561: '病' // U+75C5 <cjk>
	0x9562: '秒' // U+79D2 <cjk>
	0x9563: '苗' // U+82D7 <cjk>
	0x9564: '錨' // U+9328 <cjk>
	0x9565: '鋲' // U+92F2 <cjk>
	0x9566: '蒜' // U+849C <cjk>
	0x9567: '蛭' // U+86ED <cjk>
	0x9568: '鰭' // U+9C2D <cjk>
	0x9569: '品' // U+54C1 <cjk>
	0x956A: '彬' // U+5F6C <cjk>
	0x956B: '斌' // U+658C <cjk>
	0x956C: '浜' // U+6D5C <cjk>
	0x956D: '瀕' // U+7015 <cjk>
	0x956E: '貧' // U+8CA7 <cjk>
	0x956F: '賓' // U+8CD3 <cjk>
	0x9570: '頻' // U+983B <cjk>
	0x9571: '敏' // U+654F <cjk>
	0x9572: '瓶' // U+74F6 <cjk>
	0x9573: '不' // U+4E0D <cjk>
	0x9574: '付' // U+4ED8 <cjk>
	0x9575: '埠' // U+57E0 <cjk>
	0x9576: '夫' // U+592B <cjk>
	0x9577: '婦' // U+5A66 <cjk>
	0x9578: '富' // U+5BCC <cjk>
	0x9579: '冨' // U+51A8 <cjk>
	0x957A: '布' // U+5E03 <cjk>
	0x957B: '府' // U+5E9C <cjk>
	0x957C: '怖' // U+6016 <cjk>
	0x957D: '扶' // U+6276 <cjk>
	0x957E: '敷' // U+6577 <cjk>
	0x9580: '斧' // U+65A7 <cjk>
	0x9581: '普' // U+666E <cjk>
	0x9582: '浮' // U+6D6E <cjk>
	0x9583: '父' // U+7236 <cjk>
	0x9584: '符' // U+7B26 <cjk>
	0x9585: '腐' // U+8150 <cjk>
	0x9586: '膚' // U+819A <cjk>
	0x9587: '芙' // U+8299 <cjk>
	0x9588: '譜' // U+8B5C <cjk>
	0x9589: '負' // U+8CA0 <cjk>
	0x958A: '賦' // U+8CE6 <cjk>
	0x958B: '赴' // U+8D74 <cjk>
	0x958C: '阜' // U+961C <cjk>
	0x958D: '附' // U+9644 <cjk>
	0x958E: '侮' // U+4FAE <cjk>
	0x958F: '撫' // U+64AB <cjk>
	0x9590: '武' // U+6B66 <cjk>
	0x9591: '舞' // U+821E <cjk>
	0x9592: '葡' // U+8461 <cjk>
	0x9593: '蕪' // U+856A <cjk>
	0x9594: '部' // U+90E8 <cjk>
	0x9595: '封' // U+5C01 <cjk>
	0x9596: '楓' // U+6953 <cjk>
	0x9597: '風' // U+98A8 <cjk>
	0x9598: '葺' // U+847A <cjk>
	0x9599: '蕗' // U+8557 <cjk>
	0x959A: '伏' // U+4F0F <cjk>
	0x959B: '副' // U+526F <cjk>
	0x959C: '復' // U+5FA9 <cjk>
	0x959D: '幅' // U+5E45 <cjk>
	0x959E: '服' // U+670D <cjk>
	0x959F: '福' // U+798F <cjk>
	0x95A0: '腹' // U+8179 <cjk>
	0x95A1: '複' // U+8907 <cjk>
	0x95A2: '覆' // U+8986 <cjk>
	0x95A3: '淵' // U+6DF5 <cjk>
	0x95A4: '弗' // U+5F17 <cjk>
	0x95A5: '払' // U+6255 <cjk>
	0x95A6: '沸' // U+6CB8 <cjk>
	0x95A7: '仏' // U+4ECF <cjk>
	0x95A8: '物' // U+7269 <cjk>
	0x95A9: '鮒' // U+9B92 <cjk>
	0x95AA: '分' // U+5206 <cjk>
	0x95AB: '吻' // U+543B <cjk>
	0x95AC: '噴' // U+5674 <cjk>
	0x95AD: '墳' // U+58B3 <cjk>
	0x95AE: '憤' // U+61A4 <cjk>
	0x95AF: '扮' // U+626E <cjk>
	0x95B0: '焚' // U+711A <cjk>
	0x95B1: '奮' // U+596E <cjk>
	0x95B2: '粉' // U+7C89 <cjk>
	0x95B3: '糞' // U+7CDE <cjk>
	0x95B4: '紛' // U+7D1B <cjk>
	0x95B5: '雰' // U+96F0 <cjk>
	0x95B6: '文' // U+6587 <cjk>
	0x95B7: '聞' // U+805E <cjk>
	0x95B8: '丙' // U+4E19 <cjk>
	0x95B9: '併' // U+4F75 <cjk>
	0x95BA: '兵' // U+5175 <cjk>
	0x95BB: '塀' // U+5840 <cjk>
	0x95BC: '幣' // U+5E63 <cjk>
	0x95BD: '平' // U+5E73 <cjk>
	0x95BE: '弊' // U+5F0A <cjk>
	0x95BF: '柄' // U+67C4 <cjk>
	0x95C0: '並' // U+4E26 <cjk>
	0x95C1: '蔽' // U+853D <cjk>
	0x95C2: '閉' // U+9589 <cjk>
	0x95C3: '陛' // U+965B <cjk>
	0x95C4: '米' // U+7C73 <cjk>
	0x95C5: '頁' // U+9801 <cjk>
	0x95C6: '僻' // U+50FB <cjk>
	0x95C7: '壁' // U+58C1 <cjk>
	0x95C8: '癖' // U+7656 <cjk>
	0x95C9: '碧' // U+78A7 <cjk>
	0x95CA: '別' // U+5225 <cjk>
	0x95CB: '瞥' // U+77A5 <cjk>
	0x95CC: '蔑' // U+8511 <cjk>
	0x95CD: '箆' // U+7B86 <cjk>
	0x95CE: '偏' // U+504F <cjk>
	0x95CF: '変' // U+5909 <cjk>
	0x95D0: '片' // U+7247 <cjk>
	0x95D1: '篇' // U+7BC7 <cjk>
	0x95D2: '編' // U+7DE8 <cjk>
	0x95D3: '辺' // U+8FBA <cjk>
	0x95D4: '返' // U+8FD4 <cjk>
	0x95D5: '遍' // U+904D <cjk>
	0x95D6: '便' // U+4FBF <cjk>
	0x95D7: '勉' // U+52C9 <cjk>
	0x95D8: '娩' // U+5A29 <cjk>
	0x95D9: '弁' // U+5F01 <cjk>
	0x95DA: '鞭' // U+97AD <cjk>
	0x95DB: '保' // U+4FDD <cjk>
	0x95DC: '舗' // U+8217 <cjk>
	0x95DD: '鋪' // U+92EA <cjk>
	0x95DE: '圃' // U+5703 <cjk>
	0x95DF: '捕' // U+6355 <cjk>
	0x95E0: '歩' // U+6B69 <cjk>
	0x95E1: '甫' // U+752B <cjk>
	0x95E2: '補' // U+88DC <cjk>
	0x95E3: '輔' // U+8F14 <cjk>
	0x95E4: '穂' // U+7A42 <cjk>
	0x95E5: '募' // U+52DF <cjk>
	0x95E6: '墓' // U+5893 <cjk>
	0x95E7: '慕' // U+6155 <cjk>
	0x95E8: '戊' // U+620A <cjk>
	0x95E9: '暮' // U+66AE <cjk>
	0x95EA: '母' // U+6BCD <cjk>
	0x95EB: '簿' // U+7C3F <cjk>
	0x95EC: '菩' // U+83E9 <cjk>
	0x95ED: '倣' // U+5023 <cjk>
	0x95EE: '俸' // U+4FF8 <cjk>
	0x95EF: '包' // U+5305 <cjk>
	0x95F0: '呆' // U+5446 <cjk>
	0x95F1: '報' // U+5831 <cjk>
	0x95F2: '奉' // U+5949 <cjk>
	0x95F3: '宝' // U+5B9D <cjk>
	0x95F4: '峰' // U+5CF0 <cjk>
	0x95F5: '峯' // U+5CEF <cjk>
	0x95F6: '崩' // U+5D29 <cjk>
	0x95F7: '庖' // U+5E96 <cjk>
	0x95F8: '抱' // U+62B1 <cjk>
	0x95F9: '捧' // U+6367 <cjk>
	0x95FA: '放' // U+653E <cjk>
	0x95FB: '方' // U+65B9 <cjk>
	0x95FC: '朋' // U+670B <cjk>
	0x9640: '法' // U+6CD5 <cjk>
	0x9641: '泡' // U+6CE1 <cjk>
	0x9642: '烹' // U+70F9 <cjk>
	0x9643: '砲' // U+7832 <cjk>
	0x9644: '縫' // U+7E2B <cjk>
	0x9645: '胞' // U+80DE <cjk>
	0x9646: '芳' // U+82B3 <cjk>
	0x9647: '萌' // U+840C <cjk>
	0x9648: '蓬' // U+84EC <cjk>
	0x9649: '蜂' // U+8702 <cjk>
	0x964A: '褒' // U+8912 <cjk>
	0x964B: '訪' // U+8A2A <cjk>
	0x964C: '豊' // U+8C4A <cjk>
	0x964D: '邦' // U+90A6 <cjk>
	0x964E: '鋒' // U+92D2 <cjk>
	0x964F: '飽' // U+98FD <cjk>
	0x9650: '鳳' // U+9CF3 <cjk>
	0x9651: '鵬' // U+9D6C <cjk>
	0x9652: '乏' // U+4E4F <cjk>
	0x9653: '亡' // U+4EA1 <cjk>
	0x9654: '傍' // U+508D <cjk>
	0x9655: '剖' // U+5256 <cjk>
	0x9656: '坊' // U+574A <cjk>
	0x9657: '妨' // U+59A8 <cjk>
	0x9658: '帽' // U+5E3D <cjk>
	0x9659: '忘' // U+5FD8 <cjk>
	0x965A: '忙' // U+5FD9 <cjk>
	0x965B: '房' // U+623F <cjk>
	0x965C: '暴' // U+66B4 <cjk>
	0x965D: '望' // U+671B <cjk>
	0x965E: '某' // U+67D0 <cjk>
	0x965F: '棒' // U+68D2 <cjk>
	0x9660: '冒' // U+5192 <cjk>
	0x9661: '紡' // U+7D21 <cjk>
	0x9662: '肪' // U+80AA <cjk>
	0x9663: '膨' // U+81A8 <cjk>
	0x9664: '謀' // U+8B00 <cjk>
	0x9665: '貌' // U+8C8C <cjk>
	0x9666: '貿' // U+8CBF <cjk>
	0x9667: '鉾' // U+927E <cjk>
	0x9668: '防' // U+9632 <cjk>
	0x9669: '吠' // U+5420 <cjk>
	0x966A: '頬' // U+982C <cjk>
	0x966B: '北' // U+5317 <cjk>
	0x966C: '僕' // U+50D5 <cjk>
	0x966D: '卜' // U+535C <cjk>
	0x966E: '墨' // U+58A8 <cjk>
	0x966F: '撲' // U+64B2 <cjk>
	0x9670: '朴' // U+6734 <cjk>
	0x9671: '牧' // U+7267 <cjk>
	0x9672: '睦' // U+7766 <cjk>
	0x9673: '穆' // U+7A46 <cjk>
	0x9674: '釦' // U+91E6 <cjk>
	0x9675: '勃' // U+52C3 <cjk>
	0x9676: '没' // U+6CA1 <cjk>
	0x9677: '殆' // U+6B86 <cjk>
	0x9678: '堀' // U+5800 <cjk>
	0x9679: '幌' // U+5E4C <cjk>
	0x967A: '奔' // U+5954 <cjk>
	0x967B: '本' // U+672C <cjk>
	0x967C: '翻' // U+7FFB <cjk>
	0x967D: '凡' // U+51E1 <cjk>
	0x967E: '盆' // U+76C6 <cjk>
	0x9680: '摩' // U+6469 <cjk>
	0x9681: '磨' // U+78E8 <cjk>
	0x9682: '魔' // U+9B54 <cjk>
	0x9683: '麻' // U+9EBB <cjk>
	0x9684: '埋' // U+57CB <cjk>
	0x9685: '妹' // U+59B9 <cjk>
	0x9686: '昧' // U+6627 <cjk>
	0x9687: '枚' // U+679A <cjk>
	0x9688: '毎' // U+6BCE <cjk>
	0x9689: '哩' // U+54E9 <cjk>
	0x968A: '槙' // U+69D9 <cjk>
	0x968B: '幕' // U+5E55 <cjk>
	0x968C: '膜' // U+819C <cjk>
	0x968D: '枕' // U+6795 <cjk>
	0x968E: '鮪' // U+9BAA <cjk>
	0x968F: '柾' // U+67FE <cjk>
	0x9690: '鱒' // U+9C52 <cjk>
	0x9691: '桝' // U+685D <cjk>
	0x9692: '亦' // U+4EA6 <cjk>
	0x9693: '俣' // U+4FE3 <cjk>
	0x9694: '又' // U+53C8 <cjk>
	0x9695: '抹' // U+62B9 <cjk>
	0x9696: '末' // U+672B <cjk>
	0x9697: '沫' // U+6CAB <cjk>
	0x9698: '迄' // U+8FC4 <cjk>
	0x9699: '侭' // U+4FAD <cjk>
	0x969A: '繭' // U+7E6D <cjk>
	0x969B: '麿' // U+9EBF <cjk>
	0x969C: '万' // U+4E07 <cjk>
	0x969D: '慢' // U+6162 <cjk>
	0x969E: '満' // U+6E80 <cjk>
	0x969F: '漫' // U+6F2B <cjk>
	0x96A0: '蔓' // U+8513 <cjk>
	0x96A1: '味' // U+5473 <cjk>
	0x96A2: '未' // U+672A <cjk>
	0x96A3: '魅' // U+9B45 <cjk>
	0x96A4: '巳' // U+5DF3 <cjk>
	0x96A5: '箕' // U+7B95 <cjk>
	0x96A6: '岬' // U+5CAC <cjk>
	0x96A7: '密' // U+5BC6 <cjk>
	0x96A8: '蜜' // U+871C <cjk>
	0x96A9: '湊' // U+6E4A <cjk>
	0x96AA: '蓑' // U+84D1 <cjk>
	0x96AB: '稔' // U+7A14 <cjk>
	0x96AC: '脈' // U+8108 <cjk>
	0x96AD: '妙' // U+5999 <cjk>
	0x96AE: '粍' // U+7C8D <cjk>
	0x96AF: '民' // U+6C11 <cjk>
	0x96B0: '眠' // U+7720 <cjk>
	0x96B1: '務' // U+52D9 <cjk>
	0x96B2: '夢' // U+5922 <cjk>
	0x96B3: '無' // U+7121 <cjk>
	0x96B4: '牟' // U+725F <cjk>
	0x96B5: '矛' // U+77DB <cjk>
	0x96B6: '霧' // U+9727 <cjk>
	0x96B7: '鵡' // U+9D61 <cjk>
	0x96B8: '椋' // U+690B <cjk>
	0x96B9: '婿' // U+5A7F <cjk>
	0x96BA: '娘' // U+5A18 <cjk>
	0x96BB: '冥' // U+51A5 <cjk>
	0x96BC: '名' // U+540D <cjk>
	0x96BD: '命' // U+547D <cjk>
	0x96BE: '明' // U+660E <cjk>
	0x96BF: '盟' // U+76DF <cjk>
	0x96C0: '迷' // U+8FF7 <cjk>
	0x96C1: '銘' // U+9298 <cjk>
	0x96C2: '鳴' // U+9CF4 <cjk>
	0x96C3: '姪' // U+59EA <cjk>
	0x96C4: '牝' // U+725D <cjk>
	0x96C5: '滅' // U+6EC5 <cjk>
	0x96C6: '免' // U+514D <cjk>
	0x96C7: '棉' // U+68C9 <cjk>
	0x96C8: '綿' // U+7DBF <cjk>
	0x96C9: '緬' // U+7DEC <cjk>
	0x96CA: '面' // U+9762 <cjk>
	0x96CB: '麺' // U+9EBA <cjk>
	0x96CC: '摸' // U+6478 <cjk>
	0x96CD: '模' // U+6A21 <cjk>
	0x96CE: '茂' // U+8302 <cjk>
	0x96CF: '妄' // U+5984 <cjk>
	0x96D0: '孟' // U+5B5F <cjk>
	0x96D1: '毛' // U+6BDB <cjk>
	0x96D2: '猛' // U+731B <cjk>
	0x96D3: '盲' // U+76F2 <cjk>
	0x96D4: '網' // U+7DB2 <cjk>
	0x96D5: '耗' // U+8017 <cjk>
	0x96D6: '蒙' // U+8499 <cjk>
	0x96D7: '儲' // U+5132 <cjk>
	0x96D8: '木' // U+6728 <cjk>
	0x96D9: '黙' // U+9ED9 <cjk>
	0x96DA: '目' // U+76EE <cjk>
	0x96DB: '杢' // U+6762 <cjk>
	0x96DC: '勿' // U+52FF <cjk>
	0x96DD: '餅' // U+9905 <cjk>
	0x96DE: '尤' // U+5C24 <cjk>
	0x96DF: '戻' // U+623B <cjk>
	0x96E0: '籾' // U+7C7E <cjk>
	0x96E1: '貰' // U+8CB0 <cjk>
	0x96E2: '問' // U+554F <cjk>
	0x96E3: '悶' // U+60B6 <cjk>
	0x96E4: '紋' // U+7D0B <cjk>
	0x96E5: '門' // U+9580 <cjk>
	0x96E6: '匁' // U+5301 <cjk>
	0x96E7: '也' // U+4E5F <cjk>
	0x96E8: '冶' // U+51B6 <cjk>
	0x96E9: '夜' // U+591C <cjk>
	0x96EA: '爺' // U+723A <cjk>
	0x96EB: '耶' // U+8036 <cjk>
	0x96EC: '野' // U+91CE <cjk>
	0x96ED: '弥' // U+5F25 <cjk>
	0x96EE: '矢' // U+77E2 <cjk>
	0x96EF: '厄' // U+5384 <cjk>
	0x96F0: '役' // U+5F79 <cjk>
	0x96F1: '約' // U+7D04 <cjk>
	0x96F2: '薬' // U+85AC <cjk>
	0x96F3: '訳' // U+8A33 <cjk>
	0x96F4: '躍' // U+8E8D <cjk>
	0x96F5: '靖' // U+9756 <cjk>
	0x96F6: '柳' // U+67F3 <cjk>
	0x96F7: '薮' // U+85AE <cjk>
	0x96F8: '鑓' // U+9453 <cjk>
	0x96F9: '愉' // U+6109 <cjk>
	0x96FA: '愈' // U+6108 <cjk>
	0x96FB: '油' // U+6CB9 <cjk>
	0x96FC: '癒' // U+7652 <cjk>
	0x9740: '諭' // U+8AED <cjk>
	0x9741: '輸' // U+8F38 <cjk>
	0x9742: '唯' // U+552F <cjk>
	0x9743: '佑' // U+4F51 <cjk>
	0x9744: '優' // U+512A <cjk>
	0x9745: '勇' // U+52C7 <cjk>
	0x9746: '友' // U+53CB <cjk>
	0x9747: '宥' // U+5BA5 <cjk>
	0x9748: '幽' // U+5E7D <cjk>
	0x9749: '悠' // U+60A0 <cjk>
	0x974A: '憂' // U+6182 <cjk>
	0x974B: '揖' // U+63D6 <cjk>
	0x974C: '有' // U+6709 <cjk>
	0x974D: '柚' // U+67DA <cjk>
	0x974E: '湧' // U+6E67 <cjk>
	0x974F: '涌' // U+6D8C <cjk>
	0x9750: '猶' // U+7336 <cjk>
	0x9751: '猷' // U+7337 <cjk>
	0x9752: '由' // U+7531 <cjk>
	0x9753: '祐' // U+7950 <cjk>
	0x9754: '裕' // U+88D5 <cjk>
	0x9755: '誘' // U+8A98 <cjk>
	0x9756: '遊' // U+904A <cjk>
	0x9757: '邑' // U+9091 <cjk>
	0x9758: '郵' // U+90F5 <cjk>
	0x9759: '雄' // U+96C4 <cjk>
	0x975A: '融' // U+878D <cjk>
	0x975B: '夕' // U+5915 <cjk>
	0x975C: '予' // U+4E88 <cjk>
	0x975D: '余' // U+4F59 <cjk>
	0x975E: '与' // U+4E0E <cjk>
	0x975F: '誉' // U+8A89 <cjk>
	0x9760: '輿' // U+8F3F <cjk>
	0x9761: '預' // U+9810 <cjk>
	0x9762: '傭' // U+50AD <cjk>
	0x9763: '幼' // U+5E7C <cjk>
	0x9764: '妖' // U+5996 <cjk>
	0x9765: '容' // U+5BB9 <cjk>
	0x9766: '庸' // U+5EB8 <cjk>
	0x9767: '揚' // U+63DA <cjk>
	0x9768: '揺' // U+63FA <cjk>
	0x9769: '擁' // U+64C1 <cjk>
	0x976A: '曜' // U+66DC <cjk>
	0x976B: '楊' // U+694A <cjk>
	0x976C: '様' // U+69D8 <cjk>
	0x976D: '洋' // U+6D0B <cjk>
	0x976E: '溶' // U+6EB6 <cjk>
	0x976F: '熔' // U+7194 <cjk>
	0x9770: '用' // U+7528 <cjk>
	0x9771: '窯' // U+7AAF <cjk>
	0x9772: '羊' // U+7F8A <cjk>
	0x9773: '耀' // U+8000 <cjk>
	0x9774: '葉' // U+8449 <cjk>
	0x9775: '蓉' // U+84C9 <cjk>
	0x9776: '要' // U+8981 <cjk>
	0x9777: '謡' // U+8B21 <cjk>
	0x9778: '踊' // U+8E0A <cjk>
	0x9779: '遥' // U+9065 <cjk>
	0x977A: '陽' // U+967D <cjk>
	0x977B: '養' // U+990A <cjk>
	0x977C: '慾' // U+617E <cjk>
	0x977D: '抑' // U+6291 <cjk>
	0x977E: '欲' // U+6B32 <cjk>
	0x9780: '沃' // U+6C83 <cjk>
	0x9781: '浴' // U+6D74 <cjk>
	0x9782: '翌' // U+7FCC <cjk>
	0x9783: '翼' // U+7FFC <cjk>
	0x9784: '淀' // U+6DC0 <cjk>
	0x9785: '羅' // U+7F85 <cjk>
	0x9786: '螺' // U+87BA <cjk>
	0x9787: '裸' // U+88F8 <cjk>
	0x9788: '来' // U+6765 <cjk>
	0x9789: '莱' // U+83B1 <cjk>
	0x978A: '頼' // U+983C <cjk>
	0x978B: '雷' // U+96F7 <cjk>
	0x978C: '洛' // U+6D1B <cjk>
	0x978D: '絡' // U+7D61 <cjk>
	0x978E: '落' // U+843D <cjk>
	0x978F: '酪' // U+916A <cjk>
	0x9790: '乱' // U+4E71 <cjk>
	0x9791: '卵' // U+5375 <cjk>
	0x9792: '嵐' // U+5D50 <cjk>
	0x9793: '欄' // U+6B04 <cjk>
	0x9794: '濫' // U+6FEB <cjk>
	0x9795: '藍' // U+85CD <cjk>
	0x9796: '蘭' // U+862D <cjk>
	0x9797: '覧' // U+89A7 <cjk>
	0x9798: '利' // U+5229 <cjk>
	0x9799: '吏' // U+540F <cjk>
	0x979A: '履' // U+5C65 <cjk>
	0x979B: '李' // U+674E <cjk>
	0x979C: '梨' // U+68A8 <cjk>
	0x979D: '理' // U+7406 <cjk>
	0x979E: '璃' // U+7483 <cjk>
	0x979F: '痢' // U+75E2 <cjk>
	0x97A0: '裏' // U+88CF <cjk>
	0x97A1: '裡' // U+88E1 <cjk>
	0x97A2: '里' // U+91CC <cjk>
	0x97A3: '離' // U+96E2 <cjk>
	0x97A4: '陸' // U+9678 <cjk>
	0x97A5: '律' // U+5F8B <cjk>
	0x97A6: '率' // U+7387 <cjk>
	0x97A7: '立' // U+7ACB <cjk>
	0x97A8: '葎' // U+844E <cjk>
	0x97A9: '掠' // U+63A0 <cjk>
	0x97AA: '略' // U+7565 <cjk>
	0x97AB: '劉' // U+5289 <cjk>
	0x97AC: '流' // U+6D41 <cjk>
	0x97AD: '溜' // U+6E9C <cjk>
	0x97AE: '琉' // U+7409 <cjk>
	0x97AF: '留' // U+7559 <cjk>
	0x97B0: '硫' // U+786B <cjk>
	0x97B1: '粒' // U+7C92 <cjk>
	0x97B2: '隆' // U+9686 <cjk>
	0x97B3: '竜' // U+7ADC <cjk>
	0x97B4: '龍' // U+9F8D <cjk>
	0x97B5: '侶' // U+4FB6 <cjk>
	0x97B6: '慮' // U+616E <cjk>
	0x97B7: '旅' // U+65C5 <cjk>
	0x97B8: '虜' // U+865C <cjk>
	0x97B9: '了' // U+4E86 <cjk>
	0x97BA: '亮' // U+4EAE <cjk>
	0x97BB: '僚' // U+50DA <cjk>
	0x97BC: '両' // U+4E21 <cjk>
	0x97BD: '凌' // U+51CC <cjk>
	0x97BE: '寮' // U+5BEE <cjk>
	0x97BF: '料' // U+6599 <cjk>
	0x97C0: '梁' // U+6881 <cjk>
	0x97C1: '涼' // U+6DBC <cjk>
	0x97C2: '猟' // U+731F <cjk>
	0x97C3: '療' // U+7642 <cjk>
	0x97C4: '瞭' // U+77AD <cjk>
	0x97C5: '稜' // U+7A1C <cjk>
	0x97C6: '糧' // U+7CE7 <cjk>
	0x97C7: '良' // U+826F <cjk>
	0x97C8: '諒' // U+8AD2 <cjk>
	0x97C9: '遼' // U+907C <cjk>
	0x97CA: '量' // U+91CF <cjk>
	0x97CB: '陵' // U+9675 <cjk>
	0x97CC: '領' // U+9818 <cjk>
	0x97CD: '力' // U+529B <cjk>
	0x97CE: '緑' // U+7DD1 <cjk>
	0x97CF: '倫' // U+502B <cjk>
	0x97D0: '厘' // U+5398 <cjk>
	0x97D1: '林' // U+6797 <cjk>
	0x97D2: '淋' // U+6DCB <cjk>
	0x97D3: '燐' // U+71D0 <cjk>
	0x97D4: '琳' // U+7433 <cjk>
	0x97D5: '臨' // U+81E8 <cjk>
	0x97D6: '輪' // U+8F2A <cjk>
	0x97D7: '隣' // U+96A3 <cjk>
	0x97D8: '鱗' // U+9C57 <cjk>
	0x97D9: '麟' // U+9E9F <cjk>
	0x97DA: '瑠' // U+7460 <cjk>
	0x97DB: '塁' // U+5841 <cjk>
	0x97DC: '涙' // U+6D99 <cjk>
	0x97DD: '累' // U+7D2F <cjk>
	0x97DE: '類' // U+985E <cjk>
	0x97DF: '令' // U+4EE4 <cjk>
	0x97E0: '伶' // U+4F36 <cjk>
	0x97E1: '例' // U+4F8B <cjk>
	0x97E2: '冷' // U+51B7 <cjk>
	0x97E3: '励' // U+52B1 <cjk>
	0x97E4: '嶺' // U+5DBA <cjk>
	0x97E5: '怜' // U+601C <cjk>
	0x97E6: '玲' // U+73B2 <cjk>
	0x97E7: '礼' // U+793C <cjk>
	0x97E8: '苓' // U+82D3 <cjk>
	0x97E9: '鈴' // U+9234 <cjk>
	0x97EA: '隷' // U+96B7 <cjk>
	0x97EB: '零' // U+96F6 <cjk>
	0x97EC: '霊' // U+970A <cjk>
	0x97ED: '麗' // U+9E97 <cjk>
	0x97EE: '齢' // U+9F62 <cjk>
	0x97EF: '暦' // U+66A6 <cjk>
	0x97F0: '歴' // U+6B74 <cjk>
	0x97F1: '列' // U+5217 <cjk>
	0x97F2: '劣' // U+52A3 <cjk>
	0x97F3: '烈' // U+70C8 <cjk>
	0x97F4: '裂' // U+88C2 <cjk>
	0x97F5: '廉' // U+5EC9 <cjk>
	0x97F6: '恋' // U+604B <cjk>
	0x97F7: '憐' // U+6190 <cjk>
	0x97F8: '漣' // U+6F23 <cjk>
	0x97F9: '煉' // U+7149 <cjk>
	0x97FA: '簾' // U+7C3E <cjk>
	0x97FB: '練' // U+7DF4 <cjk>
	0x97FC: '聯' // U+806F <cjk>
	0x9840: '蓮' // U+84EE <cjk>
	0x9841: '連' // U+9023 <cjk>
	0x9842: '錬' // U+932C <cjk>
	0x9843: '呂' // U+5442 <cjk>
	0x9844: '魯' // U+9B6F <cjk>
	0x9845: '櫓' // U+6AD3 <cjk>
	0x9846: '炉' // U+7089 <cjk>
	0x9847: '賂' // U+8CC2 <cjk>
	0x9848: '路' // U+8DEF <cjk>
	0x9849: '露' // U+9732 <cjk>
	0x984A: '労' // U+52B4 <cjk>
	0x984B: '婁' // U+5A41 <cjk>
	0x984C: '廊' // U+5ECA <cjk>
	0x984D: '弄' // U+5F04 <cjk>
	0x984E: '朗' // U+6717 <cjk>
	0x984F: '楼' // U+697C <cjk>
	0x9850: '榔' // U+6994 <cjk>
	0x9851: '浪' // U+6D6A <cjk>
	0x9852: '漏' // U+6F0F <cjk>
	0x9853: '牢' // U+7262 <cjk>
	0x9854: '狼' // U+72FC <cjk>
	0x9855: '篭' // U+7BED <cjk>
	0x9856: '老' // U+8001 <cjk>
	0x9857: '聾' // U+807E <cjk>
	0x9858: '蝋' // U+874B <cjk>
	0x9859: '郎' // U+90CE <cjk>
	0x985A: '六' // U+516D <cjk>
	0x985B: '麓' // U+9E93 <cjk>
	0x985C: '禄' // U+7984 <cjk>
	0x985D: '肋' // U+808B <cjk>
	0x985E: '録' // U+9332 <cjk>
	0x985F: '論' // U+8AD6 <cjk>
	0x9860: '倭' // U+502D <cjk>
	0x9861: '和' // U+548C <cjk>
	0x9862: '話' // U+8A71 <cjk>
	0x9863: '歪' // U+6B6A <cjk>
	0x9864: '賄' // U+8CC4 <cjk>
	0x9865: '脇' // U+8107 <cjk>
	0x9866: '惑' // U+60D1 <cjk>
	0x9867: '枠' // U+67A0 <cjk>
	0x9868: '鷲' // U+9DF2 <cjk>
	0x9869: '亙' // U+4E99 <cjk>
	0x986A: '亘' // U+4E98 <cjk>
	0x986B: '鰐' // U+9C10 <cjk>
	0x986C: '詫' // U+8A6B <cjk>
	0x986D: '藁' // U+85C1 <cjk>
	0x986E: '蕨' // U+8568 <cjk>
	0x986F: '椀' // U+6900 <cjk>
	0x9870: '湾' // U+6E7E <cjk>
	0x9871: '碗' // U+7897 <cjk>
	0x9872: '腕' // U+8155 <cjk>
	0x9873: '𠮟' // U+20B9F <cjk>
	0x9874: '孁' // U+5B41 <cjk>
	0x9875: '孖' // U+5B56 <cjk>
	0x9876: '孽' // U+5B7D <cjk>
	0x9877: '宓' // U+5B93 <cjk>
	0x9878: '寘' // U+5BD8 <cjk>
	0x9879: '寬' // U+5BEC <cjk>
	0x987A: '尒' // U+5C12 <cjk>
	0x987B: '尞' // U+5C1E <cjk>
	0x987C: '尣' // U+5C23 <cjk>
	0x987D: '尫' // U+5C2B <cjk>
	0x987E: '㞍' // U+378D <cjk>
	0x9880: '屢' // U+5C62 <cjk>
	0x9881: '層' // U+FA3B CJK COMPATIBILITY IDEOGRAPH-FA3B
	0x9882: '屮' // U+FA3C CJK COMPATIBILITY IDEOGRAPH-FA3C
	0x9883: '𡚴' // U+216B4 <cjk>
	0x9884: '屺' // U+5C7A <cjk>
	0x9885: '岏' // U+5C8F <cjk>
	0x9886: '岟' // U+5C9F <cjk>
	0x9887: '岣' // U+5CA3 <cjk>
	0x9888: '岪' // U+5CAA <cjk>
	0x9889: '岺' // U+5CBA <cjk>
	0x988A: '峋' // U+5CCB <cjk>
	0x988B: '峐' // U+5CD0 <cjk>
	0x988C: '峒' // U+5CD2 <cjk>
	0x988D: '峴' // U+5CF4 <cjk>
	0x988E: '𡸴' // U+21E34 <cjk>
	0x988F: '㟢' // U+37E2 <cjk>
	0x9890: '崍' // U+5D0D <cjk>
	0x9891: '崧' // U+5D27 <cjk>
	0x9892: '﨑' // U+FA11 CJK COMPATIBILITY IDEOGRAPH-FA11
	0x9893: '嵆' // U+5D46 <cjk>
	0x9894: '嵇' // U+5D47 <cjk>
	0x9895: '嵓' // U+5D53 <cjk>
	0x9896: '嵊' // U+5D4A <cjk>
	0x9897: '嵭' // U+5D6D <cjk>
	0x9898: '嶁' // U+5D81 <cjk>
	0x9899: '嶠' // U+5DA0 <cjk>
	0x989A: '嶤' // U+5DA4 <cjk>
	0x989B: '嶧' // U+5DA7 <cjk>
	0x989C: '嶸' // U+5DB8 <cjk>
	0x989D: '巋' // U+5DCB <cjk>
	0x989E: '吞' // U+541E <cjk>
	0x989F: '弌' // U+5F0C <cjk>
	0x98A0: '丐' // U+4E10 <cjk>
	0x98A1: '丕' // U+4E15 <cjk>
	0x98A2: '个' // U+4E2A <cjk>
	0x98A3: '丱' // U+4E31 <cjk>
	0x98A4: '丶' // U+4E36 <cjk>
	0x98A5: '丼' // U+4E3C <cjk>
	0x98A6: '丿' // U+4E3F <cjk>
	0x98A7: '乂' // U+4E42 <cjk>
	0x98A8: '乖' // U+4E56 <cjk>
	0x98A9: '乘' // U+4E58 <cjk>
	0x98AA: '亂' // U+4E82 <cjk>
	0x98AB: '亅' // U+4E85 <cjk>
	0x98AC: '豫' // U+8C6B <cjk>
	0x98AD: '亊' // U+4E8A <cjk>
	0x98AE: '舒' // U+8212 <cjk>
	0x98AF: '弍' // U+5F0D <cjk>
	0x98B0: '于' // U+4E8E <cjk>
	0x98B1: '亞' // U+4E9E <cjk>
	0x98B2: '亟' // U+4E9F <cjk>
	0x98B3: '亠' // U+4EA0 <cjk>
	0x98B4: '亢' // U+4EA2 <cjk>
	0x98B5: '亰' // U+4EB0 <cjk>
	0x98B6: '亳' // U+4EB3 <cjk>
	0x98B7: '亶' // U+4EB6 <cjk>
	0x98B8: '从' // U+4ECE <cjk>
	0x98B9: '仍' // U+4ECD <cjk>
	0x98BA: '仄' // U+4EC4 <cjk>
	0x98BB: '仆' // U+4EC6 <cjk>
	0x98BC: '仂' // U+4EC2 <cjk>
	0x98BD: '仗' // U+4ED7 <cjk>
	0x98BE: '仞' // U+4EDE <cjk>
	0x98BF: '仭' // U+4EED <cjk>
	0x98C0: '仟' // U+4EDF <cjk>
	0x98C1: '价' // U+4EF7 <cjk>
	0x98C2: '伉' // U+4F09 <cjk>
	0x98C3: '佚' // U+4F5A <cjk>
	0x98C4: '估' // U+4F30 <cjk>
	0x98C5: '佛' // U+4F5B <cjk>
	0x98C6: '佝' // U+4F5D <cjk>
	0x98C7: '佗' // U+4F57 <cjk>
	0x98C8: '佇' // U+4F47 <cjk>
	0x98C9: '佶' // U+4F76 <cjk>
	0x98CA: '侈' // U+4F88 <cjk>
	0x98CB: '侏' // U+4F8F <cjk>
	0x98CC: '侘' // U+4F98 <cjk>
	0x98CD: '佻' // U+4F7B <cjk>
	0x98CE: '佩' // U+4F69 <cjk>
	0x98CF: '佰' // U+4F70 <cjk>
	0x98D0: '侑' // U+4F91 <cjk>
	0x98D1: '佯' // U+4F6F <cjk>
	0x98D2: '來' // U+4F86 <cjk>
	0x98D3: '侖' // U+4F96 <cjk>
	0x98D4: '儘' // U+5118 <cjk>
	0x98D5: '俔' // U+4FD4 <cjk>
	0x98D6: '俟' // U+4FDF <cjk>
	0x98D7: '俎' // U+4FCE <cjk>
	0x98D8: '俘' // U+4FD8 <cjk>
	0x98D9: '俛' // U+4FDB <cjk>
	0x98DA: '俑' // U+4FD1 <cjk>
	0x98DB: '俚' // U+4FDA <cjk>
	0x98DC: '俐' // U+4FD0 <cjk>
	0x98DD: '俤' // U+4FE4 <cjk>
	0x98DE: '俥' // U+4FE5 <cjk>
	0x98DF: '倚' // U+501A <cjk>
	0x98E0: '倨' // U+5028 <cjk>
	0x98E1: '倔' // U+5014 <cjk>
	0x98E2: '倪' // U+502A <cjk>
	0x98E3: '倥' // U+5025 <cjk>
	0x98E4: '倅' // U+5005 <cjk>
	0x98E5: '伜' // U+4F1C <cjk>
	0x98E6: '俶' // U+4FF6 <cjk>
	0x98E7: '倡' // U+5021 <cjk>
	0x98E8: '倩' // U+5029 <cjk>
	0x98E9: '倬' // U+502C <cjk>
	0x98EA: '俾' // U+4FFE <cjk>
	0x98EB: '俯' // U+4FEF <cjk>
	0x98EC: '們' // U+5011 <cjk>
	0x98ED: '倆' // U+5006 <cjk>
	0x98EE: '偃' // U+5043 <cjk>
	0x98EF: '假' // U+5047 <cjk>
	0x98F0: '會' // U+6703 <cjk>
	0x98F1: '偕' // U+5055 <cjk>
	0x98F2: '偐' // U+5050 <cjk>
	0x98F3: '偈' // U+5048 <cjk>
	0x98F4: '做' // U+505A <cjk>
	0x98F5: '偖' // U+5056 <cjk>
	0x98F6: '偬' // U+506C <cjk>
	0x98F7: '偸' // U+5078 <cjk>
	0x98F8: '傀' // U+5080 <cjk>
	0x98F9: '傚' // U+509A <cjk>
	0x98FA: '傅' // U+5085 <cjk>
	0x98FB: '傴' // U+50B4 <cjk>
	0x98FC: '傲' // U+50B2 <cjk>
	0x9940: '僉' // U+50C9 <cjk>
	0x9941: '僊' // U+50CA <cjk>
	0x9942: '傳' // U+50B3 <cjk>
	0x9943: '僂' // U+50C2 <cjk>
	0x9944: '僖' // U+50D6 <cjk>
	0x9945: '僞' // U+50DE <cjk>
	0x9946: '僥' // U+50E5 <cjk>
	0x9947: '僭' // U+50ED <cjk>
	0x9948: '僣' // U+50E3 <cjk>
	0x9949: '僮' // U+50EE <cjk>
	0x994A: '價' // U+50F9 <cjk>
	0x994B: '僵' // U+50F5 <cjk>
	0x994C: '儉' // U+5109 <cjk>
	0x994D: '儁' // U+5101 <cjk>
	0x994E: '儂' // U+5102 <cjk>
	0x994F: '儖' // U+5116 <cjk>
	0x9950: '儕' // U+5115 <cjk>
	0x9951: '儔' // U+5114 <cjk>
	0x9952: '儚' // U+511A <cjk>
	0x9953: '儡' // U+5121 <cjk>
	0x9954: '儺' // U+513A <cjk>
	0x9955: '儷' // U+5137 <cjk>
	0x9956: '儼' // U+513C <cjk>
	0x9957: '儻' // U+513B <cjk>
	0x9958: '儿' // U+513F <cjk>
	0x9959: '兀' // U+5140 <cjk>
	0x995A: '兒' // U+5152 <cjk>
	0x995B: '兌' // U+514C <cjk>
	0x995C: '兔' // U+5154 <cjk>
	0x995D: '兢' // U+5162 <cjk>
	0x995E: '竸' // U+7AF8 <cjk>
	0x995F: '兩' // U+5169 <cjk>
	0x9960: '兪' // U+516A <cjk>
	0x9961: '兮' // U+516E <cjk>
	0x9962: '冀' // U+5180 <cjk>
	0x9963: '冂' // U+5182 <cjk>
	0x9964: '囘' // U+56D8 <cjk>
	0x9965: '册' // U+518C <cjk>
	0x9966: '冉' // U+5189 <cjk>
	0x9967: '冏' // U+518F <cjk>
	0x9968: '冑' // U+5191 <cjk>
	0x9969: '冓' // U+5193 <cjk>
	0x996A: '冕' // U+5195 <cjk>
	0x996B: '冖' // U+5196 <cjk>
	0x996C: '冤' // U+51A4 <cjk>
	0x996D: '冦' // U+51A6 <cjk>
	0x996E: '冢' // U+51A2 <cjk>
	0x996F: '冩' // U+51A9 <cjk>
	0x9970: '冪' // U+51AA <cjk>
	0x9971: '冫' // U+51AB <cjk>
	0x9972: '决' // U+51B3 <cjk>
	0x9973: '冱' // U+51B1 <cjk>
	0x9974: '冲' // U+51B2 <cjk>
	0x9975: '冰' // U+51B0 <cjk>
	0x9976: '况' // U+51B5 <cjk>
	0x9977: '冽' // U+51BD <cjk>
	0x9978: '凅' // U+51C5 <cjk>
	0x9979: '凉' // U+51C9 <cjk>
	0x997A: '凛' // U+51DB <cjk>
	0x997B: '几' // U+51E0 <cjk>
	0x997C: '處' // U+8655 <cjk>
	0x997D: '凩' // U+51E9 <cjk>
	0x997E: '凭' // U+51ED <cjk>
	0x9980: '凰' // U+51F0 <cjk>
	0x9981: '凵' // U+51F5 <cjk>
	0x9982: '凾' // U+51FE <cjk>
	0x9983: '刄' // U+5204 <cjk>
	0x9984: '刋' // U+520B <cjk>
	0x9985: '刔' // U+5214 <cjk>
	0x9986: '刎' // U+520E <cjk>
	0x9987: '刧' // U+5227 <cjk>
	0x9988: '刪' // U+522A <cjk>
	0x9989: '刮' // U+522E <cjk>
	0x998A: '刳' // U+5233 <cjk>
	0x998B: '刹' // U+5239 <cjk>
	0x998C: '剏' // U+524F <cjk>
	0x998D: '剄' // U+5244 <cjk>
	0x998E: '剋' // U+524B <cjk>
	0x998F: '剌' // U+524C <cjk>
	0x9990: '剞' // U+525E <cjk>
	0x9991: '剔' // U+5254 <cjk>
	0x9992: '剪' // U+526A <cjk>
	0x9993: '剴' // U+5274 <cjk>
	0x9994: '剩' // U+5269 <cjk>
	0x9995: '剳' // U+5273 <cjk>
	0x9996: '剿' // U+527F <cjk>
	0x9997: '剽' // U+527D <cjk>
	0x9998: '劍' // U+528D <cjk>
	0x9999: '劔' // U+5294 <cjk>
	0x999A: '劒' // U+5292 <cjk>
	0x999B: '剱' // U+5271 <cjk>
	0x999C: '劈' // U+5288 <cjk>
	0x999D: '劑' // U+5291 <cjk>
	0x999E: '辨' // U+8FA8 <cjk>
	0x999F: '辧' // U+8FA7 <cjk>
	0x99A0: '劬' // U+52AC <cjk>
	0x99A1: '劭' // U+52AD <cjk>
	0x99A2: '劼' // U+52BC <cjk>
	0x99A3: '劵' // U+52B5 <cjk>
	0x99A4: '勁' // U+52C1 <cjk>
	0x99A5: '勍' // U+52CD <cjk>
	0x99A6: '勗' // U+52D7 <cjk>
	0x99A7: '勞' // U+52DE <cjk>
	0x99A8: '勣' // U+52E3 <cjk>
	0x99A9: '勦' // U+52E6 <cjk>
	0x99AA: '飭' // U+98ED <cjk>
	0x99AB: '勠' // U+52E0 <cjk>
	0x99AC: '勳' // U+52F3 <cjk>
	0x99AD: '勵' // U+52F5 <cjk>
	0x99AE: '勸' // U+52F8 <cjk>
	0x99AF: '勹' // U+52F9 <cjk>
	0x99B0: '匆' // U+5306 <cjk>
	0x99B1: '匈' // U+5308 <cjk>
	0x99B2: '甸' // U+7538 <cjk>
	0x99B3: '匍' // U+530D <cjk>
	0x99B4: '匐' // U+5310 <cjk>
	0x99B5: '匏' // U+530F <cjk>
	0x99B6: '匕' // U+5315 <cjk>
	0x99B7: '匚' // U+531A <cjk>
	0x99B8: '匣' // U+5323 <cjk>
	0x99B9: '匯' // U+532F <cjk>
	0x99BA: '匱' // U+5331 <cjk>
	0x99BB: '匳' // U+5333 <cjk>
	0x99BC: '匸' // U+5338 <cjk>
	0x99BD: '區' // U+5340 <cjk>
	0x99BE: '卆' // U+5346 <cjk>
	0x99BF: '卅' // U+5345 <cjk>
	0x99C0: '丗' // U+4E17 <cjk>
	0x99C1: '卉' // U+5349 <cjk>
	0x99C2: '卍' // U+534D <cjk>
	0x99C3: '凖' // U+51D6 <cjk>
	0x99C4: '卞' // U+535E <cjk>
	0x99C5: '卩' // U+5369 <cjk>
	0x99C6: '卮' // U+536E <cjk>
	0x99C7: '夘' // U+5918 <cjk>
	0x99C8: '卻' // U+537B <cjk>
	0x99C9: '卷' // U+5377 <cjk>
	0x99CA: '厂' // U+5382 <cjk>
	0x99CB: '厖' // U+5396 <cjk>
	0x99CC: '厠' // U+53A0 <cjk>
	0x99CD: '厦' // U+53A6 <cjk>
	0x99CE: '厥' // U+53A5 <cjk>
	0x99CF: '厮' // U+53AE <cjk>
	0x99D0: '厰' // U+53B0 <cjk>
	0x99D1: '厶' // U+53B6 <cjk>
	0x99D2: '參' // U+53C3 <cjk>
	0x99D3: '簒' // U+7C12 <cjk>
	0x99D4: '雙' // U+96D9 <cjk>
	0x99D5: '叟' // U+53DF <cjk>
	0x99D6: '曼' // U+66FC <cjk>
	0x99D7: '燮' // U+71EE <cjk>
	0x99D8: '叮' // U+53EE <cjk>
	0x99D9: '叨' // U+53E8 <cjk>
	0x99DA: '叭' // U+53ED <cjk>
	0x99DB: '叺' // U+53FA <cjk>
	0x99DC: '吁' // U+5401 <cjk>
	0x99DD: '吽' // U+543D <cjk>
	0x99DE: '呀' // U+5440 <cjk>
	0x99DF: '听' // U+542C <cjk>
	0x99E0: '吭' // U+542D <cjk>
	0x99E1: '吼' // U+543C <cjk>
	0x99E2: '吮' // U+542E <cjk>
	0x99E3: '吶' // U+5436 <cjk>
	0x99E4: '吩' // U+5429 <cjk>
	0x99E5: '吝' // U+541D <cjk>
	0x99E6: '呎' // U+544E <cjk>
	0x99E7: '咏' // U+548F <cjk>
	0x99E8: '呵' // U+5475 <cjk>
	0x99E9: '咎' // U+548E <cjk>
	0x99EA: '呟' // U+545F <cjk>
	0x99EB: '呱' // U+5471 <cjk>
	0x99EC: '呷' // U+5477 <cjk>
	0x99ED: '呰' // U+5470 <cjk>
	0x99EE: '咒' // U+5492 <cjk>
	0x99EF: '呻' // U+547B <cjk>
	0x99F0: '咀' // U+5480 <cjk>
	0x99F1: '呶' // U+5476 <cjk>
	0x99F2: '咄' // U+5484 <cjk>
	0x99F3: '咐' // U+5490 <cjk>
	0x99F4: '咆' // U+5486 <cjk>
	0x99F5: '哇' // U+54C7 <cjk>
	0x99F6: '咢' // U+54A2 <cjk>
	0x99F7: '咸' // U+54B8 <cjk>
	0x99F8: '咥' // U+54A5 <cjk>
	0x99F9: '咬' // U+54AC <cjk>
	0x99FA: '哄' // U+54C4 <cjk>
	0x99FB: '哈' // U+54C8 <cjk>
	0x99FC: '咨' // U+54A8 <cjk>
	0x9A40: '咫' // U+54AB <cjk>
	0x9A41: '哂' // U+54C2 <cjk>
	0x9A42: '咤' // U+54A4 <cjk>
	0x9A43: '咾' // U+54BE <cjk>
	0x9A44: '咼' // U+54BC <cjk>
	0x9A45: '哘' // U+54D8 <cjk>
	0x9A46: '哥' // U+54E5 <cjk>
	0x9A47: '哦' // U+54E6 <cjk>
	0x9A48: '唏' // U+550F <cjk>
	0x9A49: '唔' // U+5514 <cjk>
	0x9A4A: '哽' // U+54FD <cjk>
	0x9A4B: '哮' // U+54EE <cjk>
	0x9A4C: '哭' // U+54ED <cjk>
	0x9A4D: '哺' // U+54FA <cjk>
	0x9A4E: '哢' // U+54E2 <cjk>
	0x9A4F: '唹' // U+5539 <cjk>
	0x9A50: '啀' // U+5540 <cjk>
	0x9A51: '啣' // U+5563 <cjk>
	0x9A52: '啌' // U+554C <cjk>
	0x9A53: '售' // U+552E <cjk>
	0x9A54: '啜' // U+555C <cjk>
	0x9A55: '啅' // U+5545 <cjk>
	0x9A56: '啖' // U+5556 <cjk>
	0x9A57: '啗' // U+5557 <cjk>
	0x9A58: '唸' // U+5538 <cjk>
	0x9A59: '唳' // U+5533 <cjk>
	0x9A5A: '啝' // U+555D <cjk>
	0x9A5B: '喙' // U+5599 <cjk>
	0x9A5C: '喀' // U+5580 <cjk>
	0x9A5D: '咯' // U+54AF <cjk>
	0x9A5E: '喊' // U+558A <cjk>
	0x9A5F: '喟' // U+559F <cjk>
	0x9A60: '啻' // U+557B <cjk>
	0x9A61: '啾' // U+557E <cjk>
	0x9A62: '喘' // U+5598 <cjk>
	0x9A63: '喞' // U+559E <cjk>
	0x9A64: '單' // U+55AE <cjk>
	0x9A65: '啼' // U+557C <cjk>
	0x9A66: '喃' // U+5583 <cjk>
	0x9A67: '喩' // U+55A9 <cjk>
	0x9A68: '喇' // U+5587 <cjk>
	0x9A69: '喨' // U+55A8 <cjk>
	0x9A6A: '嗚' // U+55DA <cjk>
	0x9A6B: '嗅' // U+55C5 <cjk>
	0x9A6C: '嗟' // U+55DF <cjk>
	0x9A6D: '嗄' // U+55C4 <cjk>
	0x9A6E: '嗜' // U+55DC <cjk>
	0x9A6F: '嗤' // U+55E4 <cjk>
	0x9A70: '嗔' // U+55D4 <cjk>
	0x9A71: '嘔' // U+5614 <cjk>
	0x9A72: '嗷' // U+55F7 <cjk>
	0x9A73: '嘖' // U+5616 <cjk>
	0x9A74: '嗾' // U+55FE <cjk>
	0x9A75: '嗽' // U+55FD <cjk>
	0x9A76: '嘛' // U+561B <cjk>
	0x9A77: '嗹' // U+55F9 <cjk>
	0x9A78: '噎' // U+564E <cjk>
	0x9A79: '噐' // U+5650 <cjk>
	0x9A7A: '營' // U+71DF <cjk>
	0x9A7B: '嘴' // U+5634 <cjk>
	0x9A7C: '嘶' // U+5636 <cjk>
	0x9A7D: '嘲' // U+5632 <cjk>
	0x9A7E: '嘸' // U+5638 <cjk>
	0x9A80: '噫' // U+566B <cjk>
	0x9A81: '噤' // U+5664 <cjk>
	0x9A82: '嘯' // U+562F <cjk>
	0x9A83: '噬' // U+566C <cjk>
	0x9A84: '噪' // U+566A <cjk>
	0x9A85: '嚆' // U+5686 <cjk>
	0x9A86: '嚀' // U+5680 <cjk>
	0x9A87: '嚊' // U+568A <cjk>
	0x9A88: '嚠' // U+56A0 <cjk>
	0x9A89: '嚔' // U+5694 <cjk>
	0x9A8A: '嚏' // U+568F <cjk>
	0x9A8B: '嚥' // U+56A5 <cjk>
	0x9A8C: '嚮' // U+56AE <cjk>
	0x9A8D: '嚶' // U+56B6 <cjk>
	0x9A8E: '嚴' // U+56B4 <cjk>
	0x9A8F: '囂' // U+56C2 <cjk>
	0x9A90: '嚼' // U+56BC <cjk>
	0x9A91: '囁' // U+56C1 <cjk>
	0x9A92: '囃' // U+56C3 <cjk>
	0x9A93: '囀' // U+56C0 <cjk>
	0x9A94: '囈' // U+56C8 <cjk>
	0x9A95: '囎' // U+56CE <cjk>
	0x9A96: '囑' // U+56D1 <cjk>
	0x9A97: '囓' // U+56D3 <cjk>
	0x9A98: '囗' // U+56D7 <cjk>
	0x9A99: '囮' // U+56EE <cjk>
	0x9A9A: '囹' // U+56F9 <cjk>
	0x9A9B: '圀' // U+5700 <cjk>
	0x9A9C: '囿' // U+56FF <cjk>
	0x9A9D: '圄' // U+5704 <cjk>
	0x9A9E: '圉' // U+5709 <cjk>
	0x9A9F: '圈' // U+5708 <cjk>
	0x9AA0: '國' // U+570B <cjk>
	0x9AA1: '圍' // U+570D <cjk>
	0x9AA2: '圓' // U+5713 <cjk>
	0x9AA3: '團' // U+5718 <cjk>
	0x9AA4: '圖' // U+5716 <cjk>
	0x9AA5: '嗇' // U+55C7 <cjk>
	0x9AA6: '圜' // U+571C <cjk>
	0x9AA7: '圦' // U+5726 <cjk>
	0x9AA8: '圷' // U+5737 <cjk>
	0x9AA9: '圸' // U+5738 <cjk>
	0x9AAA: '坎' // U+574E <cjk>
	0x9AAB: '圻' // U+573B <cjk>
	0x9AAC: '址' // U+5740 <cjk>
	0x9AAD: '坏' // U+574F <cjk>
	0x9AAE: '坩' // U+5769 <cjk>
	0x9AAF: '埀' // U+57C0 <cjk>
	0x9AB0: '垈' // U+5788 <cjk>
	0x9AB1: '坡' // U+5761 <cjk>
	0x9AB2: '坿' // U+577F <cjk>
	0x9AB3: '垉' // U+5789 <cjk>
	0x9AB4: '垓' // U+5793 <cjk>
	0x9AB5: '垠' // U+57A0 <cjk>
	0x9AB6: '垳' // U+57B3 <cjk>
	0x9AB7: '垤' // U+57A4 <cjk>
	0x9AB8: '垪' // U+57AA <cjk>
	0x9AB9: '垰' // U+57B0 <cjk>
	0x9ABA: '埃' // U+57C3 <cjk>
	0x9ABB: '埆' // U+57C6 <cjk>
	0x9ABC: '埔' // U+57D4 <cjk>
	0x9ABD: '埒' // U+57D2 <cjk>
	0x9ABE: '埓' // U+57D3 <cjk>
	0x9ABF: '堊' // U+580A <cjk>
	0x9AC0: '埖' // U+57D6 <cjk>
	0x9AC1: '埣' // U+57E3 <cjk>
	0x9AC2: '堋' // U+580B <cjk>
	0x9AC3: '堙' // U+5819 <cjk>
	0x9AC4: '堝' // U+581D <cjk>
	0x9AC5: '塲' // U+5872 <cjk>
	0x9AC6: '堡' // U+5821 <cjk>
	0x9AC7: '塢' // U+5862 <cjk>
	0x9AC8: '塋' // U+584B <cjk>
	0x9AC9: '塰' // U+5870 <cjk>
	0x9ACA: '毀' // U+6BC0 <cjk>
	0x9ACB: '塒' // U+5852 <cjk>
	0x9ACC: '堽' // U+583D <cjk>
	0x9ACD: '塹' // U+5879 <cjk>
	0x9ACE: '墅' // U+5885 <cjk>
	0x9ACF: '墹' // U+58B9 <cjk>
	0x9AD0: '墟' // U+589F <cjk>
	0x9AD1: '墫' // U+58AB <cjk>
	0x9AD2: '墺' // U+58BA <cjk>
	0x9AD3: '壞' // U+58DE <cjk>
	0x9AD4: '墻' // U+58BB <cjk>
	0x9AD5: '墸' // U+58B8 <cjk>
	0x9AD6: '墮' // U+58AE <cjk>
	0x9AD7: '壅' // U+58C5 <cjk>
	0x9AD8: '壓' // U+58D3 <cjk>
	0x9AD9: '壑' // U+58D1 <cjk>
	0x9ADA: '壗' // U+58D7 <cjk>
	0x9ADB: '壙' // U+58D9 <cjk>
	0x9ADC: '壘' // U+58D8 <cjk>
	0x9ADD: '壥' // U+58E5 <cjk>
	0x9ADE: '壜' // U+58DC <cjk>
	0x9ADF: '壤' // U+58E4 <cjk>
	0x9AE0: '壟' // U+58DF <cjk>
	0x9AE1: '壯' // U+58EF <cjk>
	0x9AE2: '壺' // U+58FA <cjk>
	0x9AE3: '壹' // U+58F9 <cjk>
	0x9AE4: '壻' // U+58FB <cjk>
	0x9AE5: '壼' // U+58FC <cjk>
	0x9AE6: '壽' // U+58FD <cjk>
	0x9AE7: '夂' // U+5902 <cjk>
	0x9AE8: '夊' // U+590A <cjk>
	0x9AE9: '夐' // U+5910 <cjk>
	0x9AEA: '夛' // U+591B <cjk>
	0x9AEB: '梦' // U+68A6 <cjk>
	0x9AEC: '夥' // U+5925 <cjk>
	0x9AED: '夬' // U+592C <cjk>
	0x9AEE: '夭' // U+592D <cjk>
	0x9AEF: '夲' // U+5932 <cjk>
	0x9AF0: '夸' // U+5938 <cjk>
	0x9AF1: '夾' // U+593E <cjk>
	0x9AF2: '竒' // U+7AD2 <cjk>
	0x9AF3: '奕' // U+5955 <cjk>
	0x9AF4: '奐' // U+5950 <cjk>
	0x9AF5: '奎' // U+594E <cjk>
	0x9AF6: '奚' // U+595A <cjk>
	0x9AF7: '奘' // U+5958 <cjk>
	0x9AF8: '奢' // U+5962 <cjk>
	0x9AF9: '奠' // U+5960 <cjk>
	0x9AFA: '奧' // U+5967 <cjk>
	0x9AFB: '奬' // U+596C <cjk>
	0x9AFC: '奩' // U+5969 <cjk>
	0x9B40: '奸' // U+5978 <cjk>
	0x9B41: '妁' // U+5981 <cjk>
	0x9B42: '妝' // U+599D <cjk>
	0x9B43: '佞' // U+4F5E <cjk>
	0x9B44: '侫' // U+4FAB <cjk>
	0x9B45: '妣' // U+59A3 <cjk>
	0x9B46: '妲' // U+59B2 <cjk>
	0x9B47: '姆' // U+59C6 <cjk>
	0x9B48: '姨' // U+59E8 <cjk>
	0x9B49: '姜' // U+59DC <cjk>
	0x9B4A: '妍' // U+598D <cjk>
	0x9B4B: '姙' // U+59D9 <cjk>
	0x9B4C: '姚' // U+59DA <cjk>
	0x9B4D: '娥' // U+5A25 <cjk>
	0x9B4E: '娟' // U+5A1F <cjk>
	0x9B4F: '娑' // U+5A11 <cjk>
	0x9B50: '娜' // U+5A1C <cjk>
	0x9B51: '娉' // U+5A09 <cjk>
	0x9B52: '娚' // U+5A1A <cjk>
	0x9B53: '婀' // U+5A40 <cjk>
	0x9B54: '婬' // U+5A6C <cjk>
	0x9B55: '婉' // U+5A49 <cjk>
	0x9B56: '娵' // U+5A35 <cjk>
	0x9B57: '娶' // U+5A36 <cjk>
	0x9B58: '婢' // U+5A62 <cjk>
	0x9B59: '婪' // U+5A6A <cjk>
	0x9B5A: '媚' // U+5A9A <cjk>
	0x9B5B: '媼' // U+5ABC <cjk>
	0x9B5C: '媾' // U+5ABE <cjk>
	0x9B5D: '嫋' // U+5ACB <cjk>
	0x9B5E: '嫂' // U+5AC2 <cjk>
	0x9B5F: '媽' // U+5ABD <cjk>
	0x9B60: '嫣' // U+5AE3 <cjk>
	0x9B61: '嫗' // U+5AD7 <cjk>
	0x9B62: '嫦' // U+5AE6 <cjk>
	0x9B63: '嫩' // U+5AE9 <cjk>
	0x9B64: '嫖' // U+5AD6 <cjk>
	0x9B65: '嫺' // U+5AFA <cjk>
	0x9B66: '嫻' // U+5AFB <cjk>
	0x9B67: '嬌' // U+5B0C <cjk>
	0x9B68: '嬋' // U+5B0B <cjk>
	0x9B69: '嬖' // U+5B16 <cjk>
	0x9B6A: '嬲' // U+5B32 <cjk>
	0x9B6B: '嫐' // U+5AD0 <cjk>
	0x9B6C: '嬪' // U+5B2A <cjk>
	0x9B6D: '嬶' // U+5B36 <cjk>
	0x9B6E: '嬾' // U+5B3E <cjk>
	0x9B6F: '孃' // U+5B43 <cjk>
	0x9B70: '孅' // U+5B45 <cjk>
	0x9B71: '孀' // U+5B40 <cjk>
	0x9B72: '孑' // U+5B51 <cjk>
	0x9B73: '孕' // U+5B55 <cjk>
	0x9B74: '孚' // U+5B5A <cjk>
	0x9B75: '孛' // U+5B5B <cjk>
	0x9B76: '孥' // U+5B65 <cjk>
	0x9B77: '孩' // U+5B69 <cjk>
	0x9B78: '孰' // U+5B70 <cjk>
	0x9B79: '孳' // U+5B73 <cjk>
	0x9B7A: '孵' // U+5B75 <cjk>
	0x9B7B: '學' // U+5B78 <cjk>
	0x9B7C: '斈' // U+6588 <cjk>
	0x9B7D: '孺' // U+5B7A <cjk>
	0x9B7E: '宀' // U+5B80 <cjk>
	0x9B80: '它' // U+5B83 <cjk>
	0x9B81: '宦' // U+5BA6 <cjk>
	0x9B82: '宸' // U+5BB8 <cjk>
	0x9B83: '寃' // U+5BC3 <cjk>
	0x9B84: '寇' // U+5BC7 <cjk>
	0x9B85: '寉' // U+5BC9 <cjk>
	0x9B86: '寔' // U+5BD4 <cjk>
	0x9B87: '寐' // U+5BD0 <cjk>
	0x9B88: '寤' // U+5BE4 <cjk>
	0x9B89: '實' // U+5BE6 <cjk>
	0x9B8A: '寢' // U+5BE2 <cjk>
	0x9B8B: '寞' // U+5BDE <cjk>
	0x9B8C: '寥' // U+5BE5 <cjk>
	0x9B8D: '寫' // U+5BEB <cjk>
	0x9B8E: '寰' // U+5BF0 <cjk>
	0x9B8F: '寶' // U+5BF6 <cjk>
	0x9B90: '寳' // U+5BF3 <cjk>
	0x9B91: '尅' // U+5C05 <cjk>
	0x9B92: '將' // U+5C07 <cjk>
	0x9B93: '專' // U+5C08 <cjk>
	0x9B94: '對' // U+5C0D <cjk>
	0x9B95: '尓' // U+5C13 <cjk>
	0x9B96: '尠' // U+5C20 <cjk>
	0x9B97: '尢' // U+5C22 <cjk>
	0x9B98: '尨' // U+5C28 <cjk>
	0x9B99: '尸' // U+5C38 <cjk>
	0x9B9A: '尹' // U+5C39 <cjk>
	0x9B9B: '屁' // U+5C41 <cjk>
	0x9B9C: '屆' // U+5C46 <cjk>
	0x9B9D: '屎' // U+5C4E <cjk>
	0x9B9E: '屓' // U+5C53 <cjk>
	0x9B9F: '屐' // U+5C50 <cjk>
	0x9BA0: '屏' // U+5C4F <cjk>
	0x9BA1: '孱' // U+5B71 <cjk>
	0x9BA2: '屬' // U+5C6C <cjk>
	0x9BA3: '屮' // U+5C6E <cjk>
	0x9BA4: '乢' // U+4E62 <cjk>
	0x9BA5: '屶' // U+5C76 <cjk>
	0x9BA6: '屹' // U+5C79 <cjk>
	0x9BA7: '岌' // U+5C8C <cjk>
	0x9BA8: '岑' // U+5C91 <cjk>
	0x9BA9: '岔' // U+5C94 <cjk>
	0x9BAA: '妛' // U+599B <cjk>
	0x9BAB: '岫' // U+5CAB <cjk>
	0x9BAC: '岻' // U+5CBB <cjk>
	0x9BAD: '岶' // U+5CB6 <cjk>
	0x9BAE: '岼' // U+5CBC <cjk>
	0x9BAF: '岷' // U+5CB7 <cjk>
	0x9BB0: '峅' // U+5CC5 <cjk>
	0x9BB1: '岾' // U+5CBE <cjk>
	0x9BB2: '峇' // U+5CC7 <cjk>
	0x9BB3: '峙' // U+5CD9 <cjk>
	0x9BB4: '峩' // U+5CE9 <cjk>
	0x9BB5: '峽' // U+5CFD <cjk>
	0x9BB6: '峺' // U+5CFA <cjk>
	0x9BB7: '峭' // U+5CED <cjk>
	0x9BB8: '嶌' // U+5D8C <cjk>
	0x9BB9: '峪' // U+5CEA <cjk>
	0x9BBA: '崋' // U+5D0B <cjk>
	0x9BBB: '崕' // U+5D15 <cjk>
	0x9BBC: '崗' // U+5D17 <cjk>
	0x9BBD: '嵜' // U+5D5C <cjk>
	0x9BBE: '崟' // U+5D1F <cjk>
	0x9BBF: '崛' // U+5D1B <cjk>
	0x9BC0: '崑' // U+5D11 <cjk>
	0x9BC1: '崔' // U+5D14 <cjk>
	0x9BC2: '崢' // U+5D22 <cjk>
	0x9BC3: '崚' // U+5D1A <cjk>
	0x9BC4: '崙' // U+5D19 <cjk>
	0x9BC5: '崘' // U+5D18 <cjk>
	0x9BC6: '嵌' // U+5D4C <cjk>
	0x9BC7: '嵒' // U+5D52 <cjk>
	0x9BC8: '嵎' // U+5D4E <cjk>
	0x9BC9: '嵋' // U+5D4B <cjk>
	0x9BCA: '嵬' // U+5D6C <cjk>
	0x9BCB: '嵳' // U+5D73 <cjk>
	0x9BCC: '嵶' // U+5D76 <cjk>
	0x9BCD: '嶇' // U+5D87 <cjk>
	0x9BCE: '嶄' // U+5D84 <cjk>
	0x9BCF: '嶂' // U+5D82 <cjk>
	0x9BD0: '嶢' // U+5DA2 <cjk>
	0x9BD1: '嶝' // U+5D9D <cjk>
	0x9BD2: '嶬' // U+5DAC <cjk>
	0x9BD3: '嶮' // U+5DAE <cjk>
	0x9BD4: '嶽' // U+5DBD <cjk>
	0x9BD5: '嶐' // U+5D90 <cjk>
	0x9BD6: '嶷' // U+5DB7 <cjk>
	0x9BD7: '嶼' // U+5DBC <cjk>
	0x9BD8: '巉' // U+5DC9 <cjk>
	0x9BD9: '巍' // U+5DCD <cjk>
	0x9BDA: '巓' // U+5DD3 <cjk>
	0x9BDB: '巒' // U+5DD2 <cjk>
	0x9BDC: '巖' // U+5DD6 <cjk>
	0x9BDD: '巛' // U+5DDB <cjk>
	0x9BDE: '巫' // U+5DEB <cjk>
	0x9BDF: '已' // U+5DF2 <cjk>
	0x9BE0: '巵' // U+5DF5 <cjk>
	0x9BE1: '帋' // U+5E0B <cjk>
	0x9BE2: '帚' // U+5E1A <cjk>
	0x9BE3: '帙' // U+5E19 <cjk>
	0x9BE4: '帑' // U+5E11 <cjk>
	0x9BE5: '帛' // U+5E1B <cjk>
	0x9BE6: '帶' // U+5E36 <cjk>
	0x9BE7: '帷' // U+5E37 <cjk>
	0x9BE8: '幄' // U+5E44 <cjk>
	0x9BE9: '幃' // U+5E43 <cjk>
	0x9BEA: '幀' // U+5E40 <cjk>
	0x9BEB: '幎' // U+5E4E <cjk>
	0x9BEC: '幗' // U+5E57 <cjk>
	0x9BED: '幔' // U+5E54 <cjk>
	0x9BEE: '幟' // U+5E5F <cjk>
	0x9BEF: '幢' // U+5E62 <cjk>
	0x9BF0: '幤' // U+5E64 <cjk>
	0x9BF1: '幇' // U+5E47 <cjk>
	0x9BF2: '幵' // U+5E75 <cjk>
	0x9BF3: '并' // U+5E76 <cjk>
	0x9BF4: '幺' // U+5E7A <cjk>
	0x9BF5: '麼' // U+9EBC <cjk>
	0x9BF6: '广' // U+5E7F <cjk>
	0x9BF7: '庠' // U+5EA0 <cjk>
	0x9BF8: '廁' // U+5EC1 <cjk>
	0x9BF9: '廂' // U+5EC2 <cjk>
	0x9BFA: '廈' // U+5EC8 <cjk>
	0x9BFB: '廐' // U+5ED0 <cjk>
	0x9BFC: '廏' // U+5ECF <cjk>
	0x9C40: '廖' // U+5ED6 <cjk>
	0x9C41: '廣' // U+5EE3 <cjk>
	0x9C42: '廝' // U+5EDD <cjk>
	0x9C43: '廚' // U+5EDA <cjk>
	0x9C44: '廛' // U+5EDB <cjk>
	0x9C45: '廢' // U+5EE2 <cjk>
	0x9C46: '廡' // U+5EE1 <cjk>
	0x9C47: '廨' // U+5EE8 <cjk>
	0x9C48: '廩' // U+5EE9 <cjk>
	0x9C49: '廬' // U+5EEC <cjk>
	0x9C4A: '廱' // U+5EF1 <cjk>
	0x9C4B: '廳' // U+5EF3 <cjk>
	0x9C4C: '廰' // U+5EF0 <cjk>
	0x9C4D: '廴' // U+5EF4 <cjk>
	0x9C4E: '廸' // U+5EF8 <cjk>
	0x9C4F: '廾' // U+5EFE <cjk>
	0x9C50: '弃' // U+5F03 <cjk>
	0x9C51: '弉' // U+5F09 <cjk>
	0x9C52: '彝' // U+5F5D <cjk>
	0x9C53: '彜' // U+5F5C <cjk>
	0x9C54: '弋' // U+5F0B <cjk>
	0x9C55: '弑' // U+5F11 <cjk>
	0x9C56: '弖' // U+5F16 <cjk>
	0x9C57: '弩' // U+5F29 <cjk>
	0x9C58: '弭' // U+5F2D <cjk>
	0x9C59: '弸' // U+5F38 <cjk>
	0x9C5A: '彁' // U+5F41 <cjk>
	0x9C5B: '彈' // U+5F48 <cjk>
	0x9C5C: '彌' // U+5F4C <cjk>
	0x9C5D: '彎' // U+5F4E <cjk>
	0x9C5E: '弯' // U+5F2F <cjk>
	0x9C5F: '彑' // U+5F51 <cjk>
	0x9C60: '彖' // U+5F56 <cjk>
	0x9C61: '彗' // U+5F57 <cjk>
	0x9C62: '彙' // U+5F59 <cjk>
	0x9C63: '彡' // U+5F61 <cjk>
	0x9C64: '彭' // U+5F6D <cjk>
	0x9C65: '彳' // U+5F73 <cjk>
	0x9C66: '彷' // U+5F77 <cjk>
	0x9C67: '徃' // U+5F83 <cjk>
	0x9C68: '徂' // U+5F82 <cjk>
	0x9C69: '彿' // U+5F7F <cjk>
	0x9C6A: '徊' // U+5F8A <cjk>
	0x9C6B: '很' // U+5F88 <cjk>
	0x9C6C: '徑' // U+5F91 <cjk>
	0x9C6D: '徇' // U+5F87 <cjk>
	0x9C6E: '從' // U+5F9E <cjk>
	0x9C6F: '徙' // U+5F99 <cjk>
	0x9C70: '徘' // U+5F98 <cjk>
	0x9C71: '徠' // U+5FA0 <cjk>
	0x9C72: '徨' // U+5FA8 <cjk>
	0x9C73: '徭' // U+5FAD <cjk>
	0x9C74: '徼' // U+5FBC <cjk>
	0x9C75: '忖' // U+5FD6 <cjk>
	0x9C76: '忻' // U+5FFB <cjk>
	0x9C77: '忤' // U+5FE4 <cjk>
	0x9C78: '忸' // U+5FF8 <cjk>
	0x9C79: '忱' // U+5FF1 <cjk>
	0x9C7A: '忝' // U+5FDD <cjk>
	0x9C7B: '悳' // U+60B3 <cjk>
	0x9C7C: '忿' // U+5FFF <cjk>
	0x9C7D: '怡' // U+6021 <cjk>
	0x9C7E: '恠' // U+6060 <cjk>
	0x9C80: '怙' // U+6019 <cjk>
	0x9C81: '怐' // U+6010 <cjk>
	0x9C82: '怩' // U+6029 <cjk>
	0x9C83: '怎' // U+600E <cjk>
	0x9C84: '怱' // U+6031 <cjk>
	0x9C85: '怛' // U+601B <cjk>
	0x9C86: '怕' // U+6015 <cjk>
	0x9C87: '怫' // U+602B <cjk>
	0x9C88: '怦' // U+6026 <cjk>
	0x9C89: '怏' // U+600F <cjk>
	0x9C8A: '怺' // U+603A <cjk>
	0x9C8B: '恚' // U+605A <cjk>
	0x9C8C: '恁' // U+6041 <cjk>
	0x9C8D: '恪' // U+606A <cjk>
	0x9C8E: '恷' // U+6077 <cjk>
	0x9C8F: '恟' // U+605F <cjk>
	0x9C90: '恊' // U+604A <cjk>
	0x9C91: '恆' // U+6046 <cjk>
	0x9C92: '恍' // U+604D <cjk>
	0x9C93: '恣' // U+6063 <cjk>
	0x9C94: '恃' // U+6043 <cjk>
	0x9C95: '恤' // U+6064 <cjk>
	0x9C96: '恂' // U+6042 <cjk>
	0x9C97: '恬' // U+606C <cjk>
	0x9C98: '恫' // U+606B <cjk>
	0x9C99: '恙' // U+6059 <cjk>
	0x9C9A: '悁' // U+6081 <cjk>
	0x9C9B: '悍' // U+608D <cjk>
	0x9C9C: '惧' // U+60E7 <cjk>
	0x9C9D: '悃' // U+6083 <cjk>
	0x9C9E: '悚' // U+609A <cjk>
	0x9C9F: '悄' // U+6084 <cjk>
	0x9CA0: '悛' // U+609B <cjk>
	0x9CA1: '悖' // U+6096 <cjk>
	0x9CA2: '悗' // U+6097 <cjk>
	0x9CA3: '悒' // U+6092 <cjk>
	0x9CA4: '悧' // U+60A7 <cjk>
	0x9CA5: '悋' // U+608B <cjk>
	0x9CA6: '惡' // U+60E1 <cjk>
	0x9CA7: '悸' // U+60B8 <cjk>
	0x9CA8: '惠' // U+60E0 <cjk>
	0x9CA9: '惓' // U+60D3 <cjk>
	0x9CAA: '悴' // U+60B4 <cjk>
	0x9CAB: '忰' // U+5FF0 <cjk>
	0x9CAC: '悽' // U+60BD <cjk>
	0x9CAD: '惆' // U+60C6 <cjk>
	0x9CAE: '悵' // U+60B5 <cjk>
	0x9CAF: '惘' // U+60D8 <cjk>
	0x9CB0: '慍' // U+614D <cjk>
	0x9CB1: '愕' // U+6115 <cjk>
	0x9CB2: '愆' // U+6106 <cjk>
	0x9CB3: '惶' // U+60F6 <cjk>
	0x9CB4: '惷' // U+60F7 <cjk>
	0x9CB5: '愀' // U+6100 <cjk>
	0x9CB6: '惴' // U+60F4 <cjk>
	0x9CB7: '惺' // U+60FA <cjk>
	0x9CB8: '愃' // U+6103 <cjk>
	0x9CB9: '愡' // U+6121 <cjk>
	0x9CBA: '惻' // U+60FB <cjk>
	0x9CBB: '惱' // U+60F1 <cjk>
	0x9CBC: '愍' // U+610D <cjk>
	0x9CBD: '愎' // U+610E <cjk>
	0x9CBE: '慇' // U+6147 <cjk>
	0x9CBF: '愾' // U+613E <cjk>
	0x9CC0: '愨' // U+6128 <cjk>
	0x9CC1: '愧' // U+6127 <cjk>
	0x9CC2: '慊' // U+614A <cjk>
	0x9CC3: '愿' // U+613F <cjk>
	0x9CC4: '愼' // U+613C <cjk>
	0x9CC5: '愬' // U+612C <cjk>
	0x9CC6: '愴' // U+6134 <cjk>
	0x9CC7: '愽' // U+613D <cjk>
	0x9CC8: '慂' // U+6142 <cjk>
	0x9CC9: '慄' // U+6144 <cjk>
	0x9CCA: '慳' // U+6173 <cjk>
	0x9CCB: '慷' // U+6177 <cjk>
	0x9CCC: '慘' // U+6158 <cjk>
	0x9CCD: '慙' // U+6159 <cjk>
	0x9CCE: '慚' // U+615A <cjk>
	0x9CCF: '慫' // U+616B <cjk>
	0x9CD0: '慴' // U+6174 <cjk>
	0x9CD1: '慯' // U+616F <cjk>
	0x9CD2: '慥' // U+6165 <cjk>
	0x9CD3: '慱' // U+6171 <cjk>
	0x9CD4: '慟' // U+615F <cjk>
	0x9CD5: '慝' // U+615D <cjk>
	0x9CD6: '慓' // U+6153 <cjk>
	0x9CD7: '慵' // U+6175 <cjk>
	0x9CD8: '憙' // U+6199 <cjk>
	0x9CD9: '憖' // U+6196 <cjk>
	0x9CDA: '憇' // U+6187 <cjk>
	0x9CDB: '憬' // U+61AC <cjk>
	0x9CDC: '憔' // U+6194 <cjk>
	0x9CDD: '憚' // U+619A <cjk>
	0x9CDE: '憊' // U+618A <cjk>
	0x9CDF: '憑' // U+6191 <cjk>
	0x9CE0: '憫' // U+61AB <cjk>
	0x9CE1: '憮' // U+61AE <cjk>
	0x9CE2: '懌' // U+61CC <cjk>
	0x9CE3: '懊' // U+61CA <cjk>
	0x9CE4: '應' // U+61C9 <cjk>
	0x9CE5: '懷' // U+61F7 <cjk>
	0x9CE6: '懈' // U+61C8 <cjk>
	0x9CE7: '懃' // U+61C3 <cjk>
	0x9CE8: '懆' // U+61C6 <cjk>
	0x9CE9: '憺' // U+61BA <cjk>
	0x9CEA: '懋' // U+61CB <cjk>
	0x9CEB: '罹' // U+7F79 <cjk>
	0x9CEC: '懍' // U+61CD <cjk>
	0x9CED: '懦' // U+61E6 <cjk>
	0x9CEE: '懣' // U+61E3 <cjk>
	0x9CEF: '懶' // U+61F6 <cjk>
	0x9CF0: '懺' // U+61FA <cjk>
	0x9CF1: '懴' // U+61F4 <cjk>
	0x9CF2: '懿' // U+61FF <cjk>
	0x9CF3: '懽' // U+61FD <cjk>
	0x9CF4: '懼' // U+61FC <cjk>
	0x9CF5: '懾' // U+61FE <cjk>
	0x9CF6: '戀' // U+6200 <cjk>
	0x9CF7: '戈' // U+6208 <cjk>
	0x9CF8: '戉' // U+6209 <cjk>
	0x9CF9: '戍' // U+620D <cjk>
	0x9CFA: '戌' // U+620C <cjk>
	0x9CFB: '戔' // U+6214 <cjk>
	0x9CFC: '戛' // U+621B <cjk>
	0x9D40: '戞' // U+621E <cjk>
	0x9D41: '戡' // U+6221 <cjk>
	0x9D42: '截' // U+622A <cjk>
	0x9D43: '戮' // U+622E <cjk>
	0x9D44: '戰' // U+6230 <cjk>
	0x9D45: '戲' // U+6232 <cjk>
	0x9D46: '戳' // U+6233 <cjk>
	0x9D47: '扁' // U+6241 <cjk>
	0x9D48: '扎' // U+624E <cjk>
	0x9D49: '扞' // U+625E <cjk>
	0x9D4A: '扣' // U+6263 <cjk>
	0x9D4B: '扛' // U+625B <cjk>
	0x9D4C: '扠' // U+6260 <cjk>
	0x9D4D: '扨' // U+6268 <cjk>
	0x9D4E: '扼' // U+627C <cjk>
	0x9D4F: '抂' // U+6282 <cjk>
	0x9D50: '抉' // U+6289 <cjk>
	0x9D51: '找' // U+627E <cjk>
	0x9D52: '抒' // U+6292 <cjk>
	0x9D53: '抓' // U+6293 <cjk>
	0x9D54: '抖' // U+6296 <cjk>
	0x9D55: '拔' // U+62D4 <cjk>
	0x9D56: '抃' // U+6283 <cjk>
	0x9D57: '抔' // U+6294 <cjk>
	0x9D58: '拗' // U+62D7 <cjk>
	0x9D59: '拑' // U+62D1 <cjk>
	0x9D5A: '抻' // U+62BB <cjk>
	0x9D5B: '拏' // U+62CF <cjk>
	0x9D5C: '拿' // U+62FF <cjk>
	0x9D5D: '拆' // U+62C6 <cjk>
	0x9D5E: '擔' // U+64D4 <cjk>
	0x9D5F: '拈' // U+62C8 <cjk>
	0x9D60: '拜' // U+62DC <cjk>
	0x9D61: '拌' // U+62CC <cjk>
	0x9D62: '拊' // U+62CA <cjk>
	0x9D63: '拂' // U+62C2 <cjk>
	0x9D64: '拇' // U+62C7 <cjk>
	0x9D65: '抛' // U+629B <cjk>
	0x9D66: '拉' // U+62C9 <cjk>
	0x9D67: '挌' // U+630C <cjk>
	0x9D68: '拮' // U+62EE <cjk>
	0x9D69: '拱' // U+62F1 <cjk>
	0x9D6A: '挧' // U+6327 <cjk>
	0x9D6B: '挂' // U+6302 <cjk>
	0x9D6C: '挈' // U+6308 <cjk>
	0x9D6D: '拯' // U+62EF <cjk>
	0x9D6E: '拵' // U+62F5 <cjk>
	0x9D6F: '捐' // U+6350 <cjk>
	0x9D70: '挾' // U+633E <cjk>
	0x9D71: '捍' // U+634D <cjk>
	0x9D72: '搜' // U+641C <cjk>
	0x9D73: '捏' // U+634F <cjk>
	0x9D74: '掖' // U+6396 <cjk>
	0x9D75: '掎' // U+638E <cjk>
	0x9D76: '掀' // U+6380 <cjk>
	0x9D77: '掫' // U+63AB <cjk>
	0x9D78: '捶' // U+6376 <cjk>
	0x9D79: '掣' // U+63A3 <cjk>
	0x9D7A: '掏' // U+638F <cjk>
	0x9D7B: '掉' // U+6389 <cjk>
	0x9D7C: '掟' // U+639F <cjk>
	0x9D7D: '掵' // U+63B5 <cjk>
	0x9D7E: '捫' // U+636B <cjk>
	0x9D80: '捩' // U+6369 <cjk>
	0x9D81: '掾' // U+63BE <cjk>
	0x9D82: '揩' // U+63E9 <cjk>
	0x9D83: '揀' // U+63C0 <cjk>
	0x9D84: '揆' // U+63C6 <cjk>
	0x9D85: '揣' // U+63E3 <cjk>
	0x9D86: '揉' // U+63C9 <cjk>
	0x9D87: '插' // U+63D2 <cjk>
	0x9D88: '揶' // U+63F6 <cjk>
	0x9D89: '揄' // U+63C4 <cjk>
	0x9D8A: '搖' // U+6416 <cjk>
	0x9D8B: '搴' // U+6434 <cjk>
	0x9D8C: '搆' // U+6406 <cjk>
	0x9D8D: '搓' // U+6413 <cjk>
	0x9D8E: '搦' // U+6426 <cjk>
	0x9D8F: '搶' // U+6436 <cjk>
	0x9D90: '攝' // U+651D <cjk>
	0x9D91: '搗' // U+6417 <cjk>
	0x9D92: '搨' // U+6428 <cjk>
	0x9D93: '搏' // U+640F <cjk>
	0x9D94: '摧' // U+6467 <cjk>
	0x9D95: '摯' // U+646F <cjk>
	0x9D96: '摶' // U+6476 <cjk>
	0x9D97: '摎' // U+644E <cjk>
	0x9D98: '攪' // U+652A <cjk>
	0x9D99: '撕' // U+6495 <cjk>
	0x9D9A: '撓' // U+6493 <cjk>
	0x9D9B: '撥' // U+64A5 <cjk>
	0x9D9C: '撩' // U+64A9 <cjk>
	0x9D9D: '撈' // U+6488 <cjk>
	0x9D9E: '撼' // U+64BC <cjk>
	0x9D9F: '據' // U+64DA <cjk>
	0x9DA0: '擒' // U+64D2 <cjk>
	0x9DA1: '擅' // U+64C5 <cjk>
	0x9DA2: '擇' // U+64C7 <cjk>
	0x9DA3: '撻' // U+64BB <cjk>
	0x9DA4: '擘' // U+64D8 <cjk>
	0x9DA5: '擂' // U+64C2 <cjk>
	0x9DA6: '擱' // U+64F1 <cjk>
	0x9DA7: '擧' // U+64E7 <cjk>
	0x9DA8: '舉' // U+8209 <cjk>
	0x9DA9: '擠' // U+64E0 <cjk>
	0x9DAA: '擡' // U+64E1 <cjk>
	0x9DAB: '抬' // U+62AC <cjk>
	0x9DAC: '擣' // U+64E3 <cjk>
	0x9DAD: '擯' // U+64EF <cjk>
	0x9DAE: '攬' // U+652C <cjk>
	0x9DAF: '擶' // U+64F6 <cjk>
	0x9DB0: '擴' // U+64F4 <cjk>
	0x9DB1: '擲' // U+64F2 <cjk>
	0x9DB2: '擺' // U+64FA <cjk>
	0x9DB3: '攀' // U+6500 <cjk>
	0x9DB4: '擽' // U+64FD <cjk>
	0x9DB5: '攘' // U+6518 <cjk>
	0x9DB6: '攜' // U+651C <cjk>
	0x9DB7: '攅' // U+6505 <cjk>
	0x9DB8: '攤' // U+6524 <cjk>
	0x9DB9: '攣' // U+6523 <cjk>
	0x9DBA: '攫' // U+652B <cjk>
	0x9DBB: '攴' // U+6534 <cjk>
	0x9DBC: '攵' // U+6535 <cjk>
	0x9DBD: '攷' // U+6537 <cjk>
	0x9DBE: '收' // U+6536 <cjk>
	0x9DBF: '攸' // U+6538 <cjk>
	0x9DC0: '畋' // U+754B <cjk>
	0x9DC1: '效' // U+6548 <cjk>
	0x9DC2: '敖' // U+6556 <cjk>
	0x9DC3: '敕' // U+6555 <cjk>
	0x9DC4: '敍' // U+654D <cjk>
	0x9DC5: '敘' // U+6558 <cjk>
	0x9DC6: '敞' // U+655E <cjk>
	0x9DC7: '敝' // U+655D <cjk>
	0x9DC8: '敲' // U+6572 <cjk>
	0x9DC9: '數' // U+6578 <cjk>
	0x9DCA: '斂' // U+6582 <cjk>
	0x9DCB: '斃' // U+6583 <cjk>
	0x9DCC: '變' // U+8B8A <cjk>
	0x9DCD: '斛' // U+659B <cjk>
	0x9DCE: '斟' // U+659F <cjk>
	0x9DCF: '斫' // U+65AB <cjk>
	0x9DD0: '斷' // U+65B7 <cjk>
	0x9DD1: '旃' // U+65C3 <cjk>
	0x9DD2: '旆' // U+65C6 <cjk>
	0x9DD3: '旁' // U+65C1 <cjk>
	0x9DD4: '旄' // U+65C4 <cjk>
	0x9DD5: '旌' // U+65CC <cjk>
	0x9DD6: '旒' // U+65D2 <cjk>
	0x9DD7: '旛' // U+65DB <cjk>
	0x9DD8: '旙' // U+65D9 <cjk>
	0x9DD9: '无' // U+65E0 <cjk>
	0x9DDA: '旡' // U+65E1 <cjk>
	0x9DDB: '旱' // U+65F1 <cjk>
	0x9DDC: '杲' // U+6772 <cjk>
	0x9DDD: '昊' // U+660A <cjk>
	0x9DDE: '昃' // U+6603 <cjk>
	0x9DDF: '旻' // U+65FB <cjk>
	0x9DE0: '杳' // U+6773 <cjk>
	0x9DE1: '昵' // U+6635 <cjk>
	0x9DE2: '昶' // U+6636 <cjk>
	0x9DE3: '昴' // U+6634 <cjk>
	0x9DE4: '昜' // U+661C <cjk>
	0x9DE5: '晏' // U+664F <cjk>
	0x9DE6: '晄' // U+6644 <cjk>
	0x9DE7: '晉' // U+6649 <cjk>
	0x9DE8: '晁' // U+6641 <cjk>
	0x9DE9: '晞' // U+665E <cjk>
	0x9DEA: '晝' // U+665D <cjk>
	0x9DEB: '晤' // U+6664 <cjk>
	0x9DEC: '晧' // U+6667 <cjk>
	0x9DED: '晨' // U+6668 <cjk>
	0x9DEE: '晟' // U+665F <cjk>
	0x9DEF: '晢' // U+6662 <cjk>
	0x9DF0: '晰' // U+6670 <cjk>
	0x9DF1: '暃' // U+6683 <cjk>
	0x9DF2: '暈' // U+6688 <cjk>
	0x9DF3: '暎' // U+668E <cjk>
	0x9DF4: '暉' // U+6689 <cjk>
	0x9DF5: '暄' // U+6684 <cjk>
	0x9DF6: '暘' // U+6698 <cjk>
	0x9DF7: '暝' // U+669D <cjk>
	0x9DF8: '曁' // U+66C1 <cjk>
	0x9DF9: '暹' // U+66B9 <cjk>
	0x9DFA: '曉' // U+66C9 <cjk>
	0x9DFB: '暾' // U+66BE <cjk>
	0x9DFC: '暼' // U+66BC <cjk>
	0x9E40: '曄' // U+66C4 <cjk>
	0x9E41: '暸' // U+66B8 <cjk>
	0x9E42: '曖' // U+66D6 <cjk>
	0x9E43: '曚' // U+66DA <cjk>
	0x9E44: '曠' // U+66E0 <cjk>
	0x9E45: '昿' // U+663F <cjk>
	0x9E46: '曦' // U+66E6 <cjk>
	0x9E47: '曩' // U+66E9 <cjk>
	0x9E48: '曰' // U+66F0 <cjk>
	0x9E49: '曵' // U+66F5 <cjk>
	0x9E4A: '曷' // U+66F7 <cjk>
	0x9E4B: '朏' // U+670F <cjk>
	0x9E4C: '朖' // U+6716 <cjk>
	0x9E4D: '朞' // U+671E <cjk>
	0x9E4E: '朦' // U+6726 <cjk>
	0x9E4F: '朧' // U+6727 <cjk>
	0x9E50: '霸' // U+9738 <cjk>
	0x9E51: '朮' // U+672E <cjk>
	0x9E52: '朿' // U+673F <cjk>
	0x9E53: '朶' // U+6736 <cjk>
	0x9E54: '杁' // U+6741 <cjk>
	0x9E55: '朸' // U+6738 <cjk>
	0x9E56: '朷' // U+6737 <cjk>
	0x9E57: '杆' // U+6746 <cjk>
	0x9E58: '杞' // U+675E <cjk>
	0x9E59: '杠' // U+6760 <cjk>
	0x9E5A: '杙' // U+6759 <cjk>
	0x9E5B: '杣' // U+6763 <cjk>
	0x9E5C: '杤' // U+6764 <cjk>
	0x9E5D: '枉' // U+6789 <cjk>
	0x9E5E: '杰' // U+6770 <cjk>
	0x9E5F: '枩' // U+67A9 <cjk>
	0x9E60: '杼' // U+677C <cjk>
	0x9E61: '杪' // U+676A <cjk>
	0x9E62: '枌' // U+678C <cjk>
	0x9E63: '枋' // U+678B <cjk>
	0x9E64: '枦' // U+67A6 <cjk>
	0x9E65: '枡' // U+67A1 <cjk>
	0x9E66: '枅' // U+6785 <cjk>
	0x9E67: '枷' // U+67B7 <cjk>
	0x9E68: '柯' // U+67EF <cjk>
	0x9E69: '枴' // U+67B4 <cjk>
	0x9E6A: '柬' // U+67EC <cjk>
	0x9E6B: '枳' // U+67B3 <cjk>
	0x9E6C: '柩' // U+67E9 <cjk>
	0x9E6D: '枸' // U+67B8 <cjk>
	0x9E6E: '柤' // U+67E4 <cjk>
	0x9E6F: '柞' // U+67DE <cjk>
	0x9E70: '柝' // U+67DD <cjk>
	0x9E71: '柢' // U+67E2 <cjk>
	0x9E72: '柮' // U+67EE <cjk>
	0x9E73: '枹' // U+67B9 <cjk>
	0x9E74: '柎' // U+67CE <cjk>
	0x9E75: '柆' // U+67C6 <cjk>
	0x9E76: '柧' // U+67E7 <cjk>
	0x9E77: '檜' // U+6A9C <cjk>
	0x9E78: '栞' // U+681E <cjk>
	0x9E79: '框' // U+6846 <cjk>
	0x9E7A: '栩' // U+6829 <cjk>
	0x9E7B: '桀' // U+6840 <cjk>
	0x9E7C: '桍' // U+684D <cjk>
	0x9E7D: '栲' // U+6832 <cjk>
	0x9E7E: '桎' // U+684E <cjk>
	0x9E80: '梳' // U+68B3 <cjk>
	0x9E81: '栫' // U+682B <cjk>
	0x9E82: '桙' // U+6859 <cjk>
	0x9E83: '档' // U+6863 <cjk>
	0x9E84: '桷' // U+6877 <cjk>
	0x9E85: '桿' // U+687F <cjk>
	0x9E86: '梟' // U+689F <cjk>
	0x9E87: '梏' // U+688F <cjk>
	0x9E88: '梭' // U+68AD <cjk>
	0x9E89: '梔' // U+6894 <cjk>
	0x9E8A: '條' // U+689D <cjk>
	0x9E8B: '梛' // U+689B <cjk>
	0x9E8C: '梃' // U+6883 <cjk>
	0x9E8D: '檮' // U+6AAE <cjk>
	0x9E8E: '梹' // U+68B9 <cjk>
	0x9E8F: '桴' // U+6874 <cjk>
	0x9E90: '梵' // U+68B5 <cjk>
	0x9E91: '梠' // U+68A0 <cjk>
	0x9E92: '梺' // U+68BA <cjk>
	0x9E93: '椏' // U+690F <cjk>
	0x9E94: '梍' // U+688D <cjk>
	0x9E95: '桾' // U+687E <cjk>
	0x9E96: '椁' // U+6901 <cjk>
	0x9E97: '棊' // U+68CA <cjk>
	0x9E98: '椈' // U+6908 <cjk>
	0x9E99: '棘' // U+68D8 <cjk>
	0x9E9A: '椢' // U+6922 <cjk>
	0x9E9B: '椦' // U+6926 <cjk>
	0x9E9C: '棡' // U+68E1 <cjk>
	0x9E9D: '椌' // U+690C <cjk>
	0x9E9E: '棍' // U+68CD <cjk>
	0x9E9F: '棔' // U+68D4 <cjk>
	0x9EA0: '棧' // U+68E7 <cjk>
	0x9EA1: '棕' // U+68D5 <cjk>
	0x9EA2: '椶' // U+6936 <cjk>
	0x9EA3: '椒' // U+6912 <cjk>
	0x9EA4: '椄' // U+6904 <cjk>
	0x9EA5: '棗' // U+68D7 <cjk>
	0x9EA6: '棣' // U+68E3 <cjk>
	0x9EA7: '椥' // U+6925 <cjk>
	0x9EA8: '棹' // U+68F9 <cjk>
	0x9EA9: '棠' // U+68E0 <cjk>
	0x9EAA: '棯' // U+68EF <cjk>
	0x9EAB: '椨' // U+6928 <cjk>
	0x9EAC: '椪' // U+692A <cjk>
	0x9EAD: '椚' // U+691A <cjk>
	0x9EAE: '椣' // U+6923 <cjk>
	0x9EAF: '椡' // U+6921 <cjk>
	0x9EB0: '棆' // U+68C6 <cjk>
	0x9EB1: '楹' // U+6979 <cjk>
	0x9EB2: '楷' // U+6977 <cjk>
	0x9EB3: '楜' // U+695C <cjk>
	0x9EB4: '楸' // U+6978 <cjk>
	0x9EB5: '楫' // U+696B <cjk>
	0x9EB6: '楔' // U+6954 <cjk>
	0x9EB7: '楾' // U+697E <cjk>
	0x9EB8: '楮' // U+696E <cjk>
	0x9EB9: '椹' // U+6939 <cjk>
	0x9EBA: '楴' // U+6974 <cjk>
	0x9EBB: '椽' // U+693D <cjk>
	0x9EBC: '楙' // U+6959 <cjk>
	0x9EBD: '椰' // U+6930 <cjk>
	0x9EBE: '楡' // U+6961 <cjk>
	0x9EBF: '楞' // U+695E <cjk>
	0x9EC0: '楝' // U+695D <cjk>
	0x9EC1: '榁' // U+6981 <cjk>
	0x9EC2: '楪' // U+696A <cjk>
	0x9EC3: '榲' // U+69B2 <cjk>
	0x9EC4: '榮' // U+69AE <cjk>
	0x9EC5: '槐' // U+69D0 <cjk>
	0x9EC6: '榿' // U+69BF <cjk>
	0x9EC7: '槁' // U+69C1 <cjk>
	0x9EC8: '槓' // U+69D3 <cjk>
	0x9EC9: '榾' // U+69BE <cjk>
	0x9ECA: '槎' // U+69CE <cjk>
	0x9ECB: '寨' // U+5BE8 <cjk>
	0x9ECC: '槊' // U+69CA <cjk>
	0x9ECD: '槝' // U+69DD <cjk>
	0x9ECE: '榻' // U+69BB <cjk>
	0x9ECF: '槃' // U+69C3 <cjk>
	0x9ED0: '榧' // U+69A7 <cjk>
	0x9ED1: '樮' // U+6A2E <cjk>
	0x9ED2: '榑' // U+6991 <cjk>
	0x9ED3: '榠' // U+69A0 <cjk>
	0x9ED4: '榜' // U+699C <cjk>
	0x9ED5: '榕' // U+6995 <cjk>
	0x9ED6: '榴' // U+69B4 <cjk>
	0x9ED7: '槞' // U+69DE <cjk>
	0x9ED8: '槨' // U+69E8 <cjk>
	0x9ED9: '樂' // U+6A02 <cjk>
	0x9EDA: '樛' // U+6A1B <cjk>
	0x9EDB: '槿' // U+69FF <cjk>
	0x9EDC: '權' // U+6B0A <cjk>
	0x9EDD: '槹' // U+69F9 <cjk>
	0x9EDE: '槲' // U+69F2 <cjk>
	0x9EDF: '槧' // U+69E7 <cjk>
	0x9EE0: '樅' // U+6A05 <cjk>
	0x9EE1: '榱' // U+69B1 <cjk>
	0x9EE2: '樞' // U+6A1E <cjk>
	0x9EE3: '槭' // U+69ED <cjk>
	0x9EE4: '樔' // U+6A14 <cjk>
	0x9EE5: '槫' // U+69EB <cjk>
	0x9EE6: '樊' // U+6A0A <cjk>
	0x9EE7: '樒' // U+6A12 <cjk>
	0x9EE8: '櫁' // U+6AC1 <cjk>
	0x9EE9: '樣' // U+6A23 <cjk>
	0x9EEA: '樓' // U+6A13 <cjk>
	0x9EEB: '橄' // U+6A44 <cjk>
	0x9EEC: '樌' // U+6A0C <cjk>
	0x9EED: '橲' // U+6A72 <cjk>
	0x9EEE: '樶' // U+6A36 <cjk>
	0x9EEF: '橸' // U+6A78 <cjk>
	0x9EF0: '橇' // U+6A47 <cjk>
	0x9EF1: '橢' // U+6A62 <cjk>
	0x9EF2: '橙' // U+6A59 <cjk>
	0x9EF3: '橦' // U+6A66 <cjk>
	0x9EF4: '橈' // U+6A48 <cjk>
	0x9EF5: '樸' // U+6A38 <cjk>
	0x9EF6: '樢' // U+6A22 <cjk>
	0x9EF7: '檐' // U+6A90 <cjk>
	0x9EF8: '檍' // U+6A8D <cjk>
	0x9EF9: '檠' // U+6AA0 <cjk>
	0x9EFA: '檄' // U+6A84 <cjk>
	0x9EFB: '檢' // U+6AA2 <cjk>
	0x9EFC: '檣' // U+6AA3 <cjk>
	0x9F40: '檗' // U+6A97 <cjk>
	0x9F41: '蘗' // U+8617 <cjk>
	0x9F42: '檻' // U+6ABB <cjk>
	0x9F43: '櫃' // U+6AC3 <cjk>
	0x9F44: '櫂' // U+6AC2 <cjk>
	0x9F45: '檸' // U+6AB8 <cjk>
	0x9F46: '檳' // U+6AB3 <cjk>
	0x9F47: '檬' // U+6AAC <cjk>
	0x9F48: '櫞' // U+6ADE <cjk>
	0x9F49: '櫑' // U+6AD1 <cjk>
	0x9F4A: '櫟' // U+6ADF <cjk>
	0x9F4B: '檪' // U+6AAA <cjk>
	0x9F4C: '櫚' // U+6ADA <cjk>
	0x9F4D: '櫪' // U+6AEA <cjk>
	0x9F4E: '櫻' // U+6AFB <cjk>
	0x9F4F: '欅' // U+6B05 <cjk>
	0x9F50: '蘖' // U+8616 <cjk>
	0x9F51: '櫺' // U+6AFA <cjk>
	0x9F52: '欒' // U+6B12 <cjk>
	0x9F53: '欖' // U+6B16 <cjk>
	0x9F54: '鬱' // U+9B31 <cjk>
	0x9F55: '欟' // U+6B1F <cjk>
	0x9F56: '欸' // U+6B38 <cjk>
	0x9F57: '欷' // U+6B37 <cjk>
	0x9F58: '盜' // U+76DC <cjk>
	0x9F59: '欹' // U+6B39 <cjk>
	0x9F5A: '飮' // U+98EE <cjk>
	0x9F5B: '歇' // U+6B47 <cjk>
	0x9F5C: '歃' // U+6B43 <cjk>
	0x9F5D: '歉' // U+6B49 <cjk>
	0x9F5E: '歐' // U+6B50 <cjk>
	0x9F5F: '歙' // U+6B59 <cjk>
	0x9F60: '歔' // U+6B54 <cjk>
	0x9F61: '歛' // U+6B5B <cjk>
	0x9F62: '歟' // U+6B5F <cjk>
	0x9F63: '歡' // U+6B61 <cjk>
	0x9F64: '歸' // U+6B78 <cjk>
	0x9F65: '歹' // U+6B79 <cjk>
	0x9F66: '歿' // U+6B7F <cjk>
	0x9F67: '殀' // U+6B80 <cjk>
	0x9F68: '殄' // U+6B84 <cjk>
	0x9F69: '殃' // U+6B83 <cjk>
	0x9F6A: '殍' // U+6B8D <cjk>
	0x9F6B: '殘' // U+6B98 <cjk>
	0x9F6C: '殕' // U+6B95 <cjk>
	0x9F6D: '殞' // U+6B9E <cjk>
	0x9F6E: '殤' // U+6BA4 <cjk>
	0x9F6F: '殪' // U+6BAA <cjk>
	0x9F70: '殫' // U+6BAB <cjk>
	0x9F71: '殯' // U+6BAF <cjk>
	0x9F72: '殲' // U+6BB2 <cjk>
	0x9F73: '殱' // U+6BB1 <cjk>
	0x9F74: '殳' // U+6BB3 <cjk>
	0x9F75: '殷' // U+6BB7 <cjk>
	0x9F76: '殼' // U+6BBC <cjk>
	0x9F77: '毆' // U+6BC6 <cjk>
	0x9F78: '毋' // U+6BCB <cjk>
	0x9F79: '毓' // U+6BD3 <cjk>
	0x9F7A: '毟' // U+6BDF <cjk>
	0x9F7B: '毬' // U+6BEC <cjk>
	0x9F7C: '毫' // U+6BEB <cjk>
	0x9F7D: '毳' // U+6BF3 <cjk>
	0x9F7E: '毯' // U+6BEF <cjk>
	0x9F80: '麾' // U+9EBE <cjk>
	0x9F81: '氈' // U+6C08 <cjk>
	0x9F82: '氓' // U+6C13 <cjk>
	0x9F83: '气' // U+6C14 <cjk>
	0x9F84: '氛' // U+6C1B <cjk>
	0x9F85: '氤' // U+6C24 <cjk>
	0x9F86: '氣' // U+6C23 <cjk>
	0x9F87: '汞' // U+6C5E <cjk>
	0x9F88: '汕' // U+6C55 <cjk>
	0x9F89: '汢' // U+6C62 <cjk>
	0x9F8A: '汪' // U+6C6A <cjk>
	0x9F8B: '沂' // U+6C82 <cjk>
	0x9F8C: '沍' // U+6C8D <cjk>
	0x9F8D: '沚' // U+6C9A <cjk>
	0x9F8E: '沁' // U+6C81 <cjk>
	0x9F8F: '沛' // U+6C9B <cjk>
	0x9F90: '汾' // U+6C7E <cjk>
	0x9F91: '汨' // U+6C68 <cjk>
	0x9F92: '汳' // U+6C73 <cjk>
	0x9F93: '沒' // U+6C92 <cjk>
	0x9F94: '沐' // U+6C90 <cjk>
	0x9F95: '泄' // U+6CC4 <cjk>
	0x9F96: '泱' // U+6CF1 <cjk>
	0x9F97: '泓' // U+6CD3 <cjk>
	0x9F98: '沽' // U+6CBD <cjk>
	0x9F99: '泗' // U+6CD7 <cjk>
	0x9F9A: '泅' // U+6CC5 <cjk>
	0x9F9B: '泝' // U+6CDD <cjk>
	0x9F9C: '沮' // U+6CAE <cjk>
	0x9F9D: '沱' // U+6CB1 <cjk>
	0x9F9E: '沾' // U+6CBE <cjk>
	0x9F9F: '沺' // U+6CBA <cjk>
	0x9FA0: '泛' // U+6CDB <cjk>
	0x9FA1: '泯' // U+6CEF <cjk>
	0x9FA2: '泙' // U+6CD9 <cjk>
	0x9FA3: '泪' // U+6CEA <cjk>
	0x9FA4: '洟' // U+6D1F <cjk>
	0x9FA5: '衍' // U+884D <cjk>
	0x9FA6: '洶' // U+6D36 <cjk>
	0x9FA7: '洫' // U+6D2B <cjk>
	0x9FA8: '洽' // U+6D3D <cjk>
	0x9FA9: '洸' // U+6D38 <cjk>
	0x9FAA: '洙' // U+6D19 <cjk>
	0x9FAB: '洵' // U+6D35 <cjk>
	0x9FAC: '洳' // U+6D33 <cjk>
	0x9FAD: '洒' // U+6D12 <cjk>
	0x9FAE: '洌' // U+6D0C <cjk>
	0x9FAF: '浣' // U+6D63 <cjk>
	0x9FB0: '涓' // U+6D93 <cjk>
	0x9FB1: '浤' // U+6D64 <cjk>
	0x9FB2: '浚' // U+6D5A <cjk>
	0x9FB3: '浹' // U+6D79 <cjk>
	0x9FB4: '浙' // U+6D59 <cjk>
	0x9FB5: '涎' // U+6D8E <cjk>
	0x9FB6: '涕' // U+6D95 <cjk>
	0x9FB7: '濤' // U+6FE4 <cjk>
	0x9FB8: '涅' // U+6D85 <cjk>
	0x9FB9: '淹' // U+6DF9 <cjk>
	0x9FBA: '渕' // U+6E15 <cjk>
	0x9FBB: '渊' // U+6E0A <cjk>
	0x9FBC: '涵' // U+6DB5 <cjk>
	0x9FBD: '淇' // U+6DC7 <cjk>
	0x9FBE: '淦' // U+6DE6 <cjk>
	0x9FBF: '涸' // U+6DB8 <cjk>
	0x9FC0: '淆' // U+6DC6 <cjk>
	0x9FC1: '淬' // U+6DEC <cjk>
	0x9FC2: '淞' // U+6DDE <cjk>
	0x9FC3: '淌' // U+6DCC <cjk>
	0x9FC4: '淨' // U+6DE8 <cjk>
	0x9FC5: '淒' // U+6DD2 <cjk>
	0x9FC6: '淅' // U+6DC5 <cjk>
	0x9FC7: '淺' // U+6DFA <cjk>
	0x9FC8: '淙' // U+6DD9 <cjk>
	0x9FC9: '淤' // U+6DE4 <cjk>
	0x9FCA: '淕' // U+6DD5 <cjk>
	0x9FCB: '淪' // U+6DEA <cjk>
	0x9FCC: '淮' // U+6DEE <cjk>
	0x9FCD: '渭' // U+6E2D <cjk>
	0x9FCE: '湮' // U+6E6E <cjk>
	0x9FCF: '渮' // U+6E2E <cjk>
	0x9FD0: '渙' // U+6E19 <cjk>
	0x9FD1: '湲' // U+6E72 <cjk>
	0x9FD2: '湟' // U+6E5F <cjk>
	0x9FD3: '渾' // U+6E3E <cjk>
	0x9FD4: '渣' // U+6E23 <cjk>
	0x9FD5: '湫' // U+6E6B <cjk>
	0x9FD6: '渫' // U+6E2B <cjk>
	0x9FD7: '湶' // U+6E76 <cjk>
	0x9FD8: '湍' // U+6E4D <cjk>
	0x9FD9: '渟' // U+6E1F <cjk>
	0x9FDA: '湃' // U+6E43 <cjk>
	0x9FDB: '渺' // U+6E3A <cjk>
	0x9FDC: '湎' // U+6E4E <cjk>
	0x9FDD: '渤' // U+6E24 <cjk>
	0x9FDE: '滿' // U+6EFF <cjk>
	0x9FDF: '渝' // U+6E1D <cjk>
	0x9FE0: '游' // U+6E38 <cjk>
	0x9FE1: '溂' // U+6E82 <cjk>
	0x9FE2: '溪' // U+6EAA <cjk>
	0x9FE3: '溘' // U+6E98 <cjk>
	0x9FE4: '滉' // U+6EC9 <cjk>
	0x9FE5: '溷' // U+6EB7 <cjk>
	0x9FE6: '滓' // U+6ED3 <cjk>
	0x9FE7: '溽' // U+6EBD <cjk>
	0x9FE8: '溯' // U+6EAF <cjk>
	0x9FE9: '滄' // U+6EC4 <cjk>
	0x9FEA: '溲' // U+6EB2 <cjk>
	0x9FEB: '滔' // U+6ED4 <cjk>
	0x9FEC: '滕' // U+6ED5 <cjk>
	0x9FED: '溏' // U+6E8F <cjk>
	0x9FEE: '溥' // U+6EA5 <cjk>
	0x9FEF: '滂' // U+6EC2 <cjk>
	0x9FF0: '溟' // U+6E9F <cjk>
	0x9FF1: '潁' // U+6F41 <cjk>
	0x9FF2: '漑' // U+6F11 <cjk>
	0x9FF3: '灌' // U+704C <cjk>
	0x9FF4: '滬' // U+6EEC <cjk>
	0x9FF5: '滸' // U+6EF8 <cjk>
	0x9FF6: '滾' // U+6EFE <cjk>
	0x9FF7: '漿' // U+6F3F <cjk>
	0x9FF8: '滲' // U+6EF2 <cjk>
	0x9FF9: '漱' // U+6F31 <cjk>
	0x9FFA: '滯' // U+6EEF <cjk>
	0x9FFB: '漲' // U+6F32 <cjk>
	0x9FFC: '滌' // U+6ECC <cjk>
	0xE040: '漾' // U+6F3E <cjk>
	0xE041: '漓' // U+6F13 <cjk>
	0xE042: '滷' // U+6EF7 <cjk>
	0xE043: '澆' // U+6F86 <cjk>
	0xE044: '潺' // U+6F7A <cjk>
	0xE045: '潸' // U+6F78 <cjk>
	0xE046: '澁' // U+6F81 <cjk>
	0xE047: '澀' // U+6F80 <cjk>
	0xE048: '潯' // U+6F6F <cjk>
	0xE049: '潛' // U+6F5B <cjk>
	0xE04A: '濳' // U+6FF3 <cjk>
	0xE04B: '潭' // U+6F6D <cjk>
	0xE04C: '澂' // U+6F82 <cjk>
	0xE04D: '潼' // U+6F7C <cjk>
	0xE04E: '潘' // U+6F58 <cjk>
	0xE04F: '澎' // U+6F8E <cjk>
	0xE050: '澑' // U+6F91 <cjk>
	0xE051: '濂' // U+6FC2 <cjk>
	0xE052: '潦' // U+6F66 <cjk>
	0xE053: '澳' // U+6FB3 <cjk>
	0xE054: '澣' // U+6FA3 <cjk>
	0xE055: '澡' // U+6FA1 <cjk>
	0xE056: '澤' // U+6FA4 <cjk>
	0xE057: '澹' // U+6FB9 <cjk>
	0xE058: '濆' // U+6FC6 <cjk>
	0xE059: '澪' // U+6FAA <cjk>
	0xE05A: '濟' // U+6FDF <cjk>
	0xE05B: '濕' // U+6FD5 <cjk>
	0xE05C: '濬' // U+6FEC <cjk>
	0xE05D: '濔' // U+6FD4 <cjk>
	0xE05E: '濘' // U+6FD8 <cjk>
	0xE05F: '濱' // U+6FF1 <cjk>
	0xE060: '濮' // U+6FEE <cjk>
	0xE061: '濛' // U+6FDB <cjk>
	0xE062: '瀉' // U+7009 <cjk>
	0xE063: '瀋' // U+700B <cjk>
	0xE064: '濺' // U+6FFA <cjk>
	0xE065: '瀑' // U+7011 <cjk>
	0xE066: '瀁' // U+7001 <cjk>
	0xE067: '瀏' // U+700F <cjk>
	0xE068: '濾' // U+6FFE <cjk>
	0xE069: '瀛' // U+701B <cjk>
	0xE06A: '瀚' // U+701A <cjk>
	0xE06B: '潴' // U+6F74 <cjk>
	0xE06C: '瀝' // U+701D <cjk>
	0xE06D: '瀘' // U+7018 <cjk>
	0xE06E: '瀟' // U+701F <cjk>
	0xE06F: '瀰' // U+7030 <cjk>
	0xE070: '瀾' // U+703E <cjk>
	0xE071: '瀲' // U+7032 <cjk>
	0xE072: '灑' // U+7051 <cjk>
	0xE073: '灣' // U+7063 <cjk>
	0xE074: '炙' // U+7099 <cjk>
	0xE075: '炒' // U+7092 <cjk>
	0xE076: '炯' // U+70AF <cjk>
	0xE077: '烱' // U+70F1 <cjk>
	0xE078: '炬' // U+70AC <cjk>
	0xE079: '炸' // U+70B8 <cjk>
	0xE07A: '炳' // U+70B3 <cjk>
	0xE07B: '炮' // U+70AE <cjk>
	0xE07C: '烟' // U+70DF <cjk>
	0xE07D: '烋' // U+70CB <cjk>
	0xE07E: '烝' // U+70DD <cjk>
	0xE080: '烙' // U+70D9 <cjk>
	0xE081: '焉' // U+7109 <cjk>
	0xE082: '烽' // U+70FD <cjk>
	0xE083: '焜' // U+711C <cjk>
	0xE084: '焙' // U+7119 <cjk>
	0xE085: '煥' // U+7165 <cjk>
	0xE086: '煕' // U+7155 <cjk>
	0xE087: '熈' // U+7188 <cjk>
	0xE088: '煦' // U+7166 <cjk>
	0xE089: '煢' // U+7162 <cjk>
	0xE08A: '煌' // U+714C <cjk>
	0xE08B: '煖' // U+7156 <cjk>
	0xE08C: '煬' // U+716C <cjk>
	0xE08D: '熏' // U+718F <cjk>
	0xE08E: '燻' // U+71FB <cjk>
	0xE08F: '熄' // U+7184 <cjk>
	0xE090: '熕' // U+7195 <cjk>
	0xE091: '熨' // U+71A8 <cjk>
	0xE092: '熬' // U+71AC <cjk>
	0xE093: '燗' // U+71D7 <cjk>
	0xE094: '熹' // U+71B9 <cjk>
	0xE095: '熾' // U+71BE <cjk>
	0xE096: '燒' // U+71D2 <cjk>
	0xE097: '燉' // U+71C9 <cjk>
	0xE098: '燔' // U+71D4 <cjk>
	0xE099: '燎' // U+71CE <cjk>
	0xE09A: '燠' // U+71E0 <cjk>
	0xE09B: '燬' // U+71EC <cjk>
	0xE09C: '燧' // U+71E7 <cjk>
	0xE09D: '燵' // U+71F5 <cjk>
	0xE09E: '燼' // U+71FC <cjk>
	0xE09F: '燹' // U+71F9 <cjk>
	0xE0A0: '燿' // U+71FF <cjk>
	0xE0A1: '爍' // U+720D <cjk>
	0xE0A2: '爐' // U+7210 <cjk>
	0xE0A3: '爛' // U+721B <cjk>
	0xE0A4: '爨' // U+7228 <cjk>
	0xE0A5: '爭' // U+722D <cjk>
	0xE0A6: '爬' // U+722C <cjk>
	0xE0A7: '爰' // U+7230 <cjk>
	0xE0A8: '爲' // U+7232 <cjk>
	0xE0A9: '爻' // U+723B <cjk>
	0xE0AA: '爼' // U+723C <cjk>
	0xE0AB: '爿' // U+723F <cjk>
	0xE0AC: '牀' // U+7240 <cjk>
	0xE0AD: '牆' // U+7246 <cjk>
	0xE0AE: '牋' // U+724B <cjk>
	0xE0AF: '牘' // U+7258 <cjk>
	0xE0B0: '牴' // U+7274 <cjk>
	0xE0B1: '牾' // U+727E <cjk>
	0xE0B2: '犂' // U+7282 <cjk>
	0xE0B3: '犁' // U+7281 <cjk>
	0xE0B4: '犇' // U+7287 <cjk>
	0xE0B5: '犒' // U+7292 <cjk>
	0xE0B6: '犖' // U+7296 <cjk>
	0xE0B7: '犢' // U+72A2 <cjk>
	0xE0B8: '犧' // U+72A7 <cjk>
	0xE0B9: '犹' // U+72B9 <cjk>
	0xE0BA: '犲' // U+72B2 <cjk>
	0xE0BB: '狃' // U+72C3 <cjk>
	0xE0BC: '狆' // U+72C6 <cjk>
	0xE0BD: '狄' // U+72C4 <cjk>
	0xE0BE: '狎' // U+72CE <cjk>
	0xE0BF: '狒' // U+72D2 <cjk>
	0xE0C0: '狢' // U+72E2 <cjk>
	0xE0C1: '狠' // U+72E0 <cjk>
	0xE0C2: '狡' // U+72E1 <cjk>
	0xE0C3: '狹' // U+72F9 <cjk>
	0xE0C4: '狷' // U+72F7 <cjk>
	0xE0C5: '倏' // U+500F <cjk>
	0xE0C6: '猗' // U+7317 <cjk>
	0xE0C7: '猊' // U+730A <cjk>
	0xE0C8: '猜' // U+731C <cjk>
	0xE0C9: '猖' // U+7316 <cjk>
	0xE0CA: '猝' // U+731D <cjk>
	0xE0CB: '猴' // U+7334 <cjk>
	0xE0CC: '猯' // U+732F <cjk>
	0xE0CD: '猩' // U+7329 <cjk>
	0xE0CE: '猥' // U+7325 <cjk>
	0xE0CF: '猾' // U+733E <cjk>
	0xE0D0: '獎' // U+734E <cjk>
	0xE0D1: '獏' // U+734F <cjk>
	0xE0D2: '默' // U+9ED8 <cjk>
	0xE0D3: '獗' // U+7357 <cjk>
	0xE0D4: '獪' // U+736A <cjk>
	0xE0D5: '獨' // U+7368 <cjk>
	0xE0D6: '獰' // U+7370 <cjk>
	0xE0D7: '獸' // U+7378 <cjk>
	0xE0D8: '獵' // U+7375 <cjk>
	0xE0D9: '獻' // U+737B <cjk>
	0xE0DA: '獺' // U+737A <cjk>
	0xE0DB: '珈' // U+73C8 <cjk>
	0xE0DC: '玳' // U+73B3 <cjk>
	0xE0DD: '珎' // U+73CE <cjk>
	0xE0DE: '玻' // U+73BB <cjk>
	0xE0DF: '珀' // U+73C0 <cjk>
	0xE0E0: '珥' // U+73E5 <cjk>
	0xE0E1: '珮' // U+73EE <cjk>
	0xE0E2: '珞' // U+73DE <cjk>
	0xE0E3: '璢' // U+74A2 <cjk>
	0xE0E4: '琅' // U+7405 <cjk>
	0xE0E5: '瑯' // U+746F <cjk>
	0xE0E6: '琥' // U+7425 <cjk>
	0xE0E7: '珸' // U+73F8 <cjk>
	0xE0E8: '琲' // U+7432 <cjk>
	0xE0E9: '琺' // U+743A <cjk>
	0xE0EA: '瑕' // U+7455 <cjk>
	0xE0EB: '琿' // U+743F <cjk>
	0xE0EC: '瑟' // U+745F <cjk>
	0xE0ED: '瑙' // U+7459 <cjk>
	0xE0EE: '瑁' // U+7441 <cjk>
	0xE0EF: '瑜' // U+745C <cjk>
	0xE0F0: '瑩' // U+7469 <cjk>
	0xE0F1: '瑰' // U+7470 <cjk>
	0xE0F2: '瑣' // U+7463 <cjk>
	0xE0F3: '瑪' // U+746A <cjk>
	0xE0F4: '瑶' // U+7476 <cjk>
	0xE0F5: '瑾' // U+747E <cjk>
	0xE0F6: '璋' // U+748B <cjk>
	0xE0F7: '璞' // U+749E <cjk>
	0xE0F8: '璧' // U+74A7 <cjk>
	0xE0F9: '瓊' // U+74CA <cjk>
	0xE0FA: '瓏' // U+74CF <cjk>
	0xE0FB: '瓔' // U+74D4 <cjk>
	0xE0FC: '珱' // U+73F1 <cjk>
	0xE140: '瓠' // U+74E0 <cjk>
	0xE141: '瓣' // U+74E3 <cjk>
	0xE142: '瓧' // U+74E7 <cjk>
	0xE143: '瓩' // U+74E9 <cjk>
	0xE144: '瓮' // U+74EE <cjk>
	0xE145: '瓲' // U+74F2 <cjk>
	0xE146: '瓰' // U+74F0 <cjk>
	0xE147: '瓱' // U+74F1 <cjk>
	0xE148: '瓸' // U+74F8 <cjk>
	0xE149: '瓷' // U+74F7 <cjk>
	0xE14A: '甄' // U+7504 <cjk>
	0xE14B: '甃' // U+7503 <cjk>
	0xE14C: '甅' // U+7505 <cjk>
	0xE14D: '甌' // U+750C <cjk>
	0xE14E: '甎' // U+750E <cjk>
	0xE14F: '甍' // U+750D <cjk>
	0xE150: '甕' // U+7515 <cjk>
	0xE151: '甓' // U+7513 <cjk>
	0xE152: '甞' // U+751E <cjk>
	0xE153: '甦' // U+7526 <cjk>
	0xE154: '甬' // U+752C <cjk>
	0xE155: '甼' // U+753C <cjk>
	0xE156: '畄' // U+7544 <cjk>
	0xE157: '畍' // U+754D <cjk>
	0xE158: '畊' // U+754A <cjk>
	0xE159: '畉' // U+7549 <cjk>
	0xE15A: '畛' // U+755B <cjk>
	0xE15B: '畆' // U+7546 <cjk>
	0xE15C: '畚' // U+755A <cjk>
	0xE15D: '畩' // U+7569 <cjk>
	0xE15E: '畤' // U+7564 <cjk>
	0xE15F: '畧' // U+7567 <cjk>
	0xE160: '畫' // U+756B <cjk>
	0xE161: '畭' // U+756D <cjk>
	0xE162: '畸' // U+7578 <cjk>
	0xE163: '當' // U+7576 <cjk>
	0xE164: '疆' // U+7586 <cjk>
	0xE165: '疇' // U+7587 <cjk>
	0xE166: '畴' // U+7574 <cjk>
	0xE167: '疊' // U+758A <cjk>
	0xE168: '疉' // U+7589 <cjk>
	0xE169: '疂' // U+7582 <cjk>
	0xE16A: '疔' // U+7594 <cjk>
	0xE16B: '疚' // U+759A <cjk>
	0xE16C: '疝' // U+759D <cjk>
	0xE16D: '疥' // U+75A5 <cjk>
	0xE16E: '疣' // U+75A3 <cjk>
	0xE16F: '痂' // U+75C2 <cjk>
	0xE170: '疳' // U+75B3 <cjk>
	0xE171: '痃' // U+75C3 <cjk>
	0xE172: '疵' // U+75B5 <cjk>
	0xE173: '疽' // U+75BD <cjk>
	0xE174: '疸' // U+75B8 <cjk>
	0xE175: '疼' // U+75BC <cjk>
	0xE176: '疱' // U+75B1 <cjk>
	0xE177: '痍' // U+75CD <cjk>
	0xE178: '痊' // U+75CA <cjk>
	0xE179: '痒' // U+75D2 <cjk>
	0xE17A: '痙' // U+75D9 <cjk>
	0xE17B: '痣' // U+75E3 <cjk>
	0xE17C: '痞' // U+75DE <cjk>
	0xE17D: '痾' // U+75FE <cjk>
	0xE17E: '痿' // U+75FF <cjk>
	0xE180: '痼' // U+75FC <cjk>
	0xE181: '瘁' // U+7601 <cjk>
	0xE182: '痰' // U+75F0 <cjk>
	0xE183: '痺' // U+75FA <cjk>
	0xE184: '痲' // U+75F2 <cjk>
	0xE185: '痳' // U+75F3 <cjk>
	0xE186: '瘋' // U+760B <cjk>
	0xE187: '瘍' // U+760D <cjk>
	0xE188: '瘉' // U+7609 <cjk>
	0xE189: '瘟' // U+761F <cjk>
	0xE18A: '瘧' // U+7627 <cjk>
	0xE18B: '瘠' // U+7620 <cjk>
	0xE18C: '瘡' // U+7621 <cjk>
	0xE18D: '瘢' // U+7622 <cjk>
	0xE18E: '瘤' // U+7624 <cjk>
	0xE18F: '瘴' // U+7634 <cjk>
	0xE190: '瘰' // U+7630 <cjk>
	0xE191: '瘻' // U+763B <cjk>
	0xE192: '癇' // U+7647 <cjk>
	0xE193: '癈' // U+7648 <cjk>
	0xE194: '癆' // U+7646 <cjk>
	0xE195: '癜' // U+765C <cjk>
	0xE196: '癘' // U+7658 <cjk>
	0xE197: '癡' // U+7661 <cjk>
	0xE198: '癢' // U+7662 <cjk>
	0xE199: '癨' // U+7668 <cjk>
	0xE19A: '癩' // U+7669 <cjk>
	0xE19B: '癪' // U+766A <cjk>
	0xE19C: '癧' // U+7667 <cjk>
	0xE19D: '癬' // U+766C <cjk>
	0xE19E: '癰' // U+7670 <cjk>
	0xE19F: '癲' // U+7672 <cjk>
	0xE1A0: '癶' // U+7676 <cjk>
	0xE1A1: '癸' // U+7678 <cjk>
	0xE1A2: '發' // U+767C <cjk>
	0xE1A3: '皀' // U+7680 <cjk>
	0xE1A4: '皃' // U+7683 <cjk>
	0xE1A5: '皈' // U+7688 <cjk>
	0xE1A6: '皋' // U+768B <cjk>
	0xE1A7: '皎' // U+768E <cjk>
	0xE1A8: '皖' // U+7696 <cjk>
	0xE1A9: '皓' // U+7693 <cjk>
	0xE1AA: '皙' // U+7699 <cjk>
	0xE1AB: '皚' // U+769A <cjk>
	0xE1AC: '皰' // U+76B0 <cjk>
	0xE1AD: '皴' // U+76B4 <cjk>
	0xE1AE: '皸' // U+76B8 <cjk>
	0xE1AF: '皹' // U+76B9 <cjk>
	0xE1B0: '皺' // U+76BA <cjk>
	0xE1B1: '盂' // U+76C2 <cjk>
	0xE1B2: '盍' // U+76CD <cjk>
	0xE1B3: '盖' // U+76D6 <cjk>
	0xE1B4: '盒' // U+76D2 <cjk>
	0xE1B5: '盞' // U+76DE <cjk>
	0xE1B6: '盡' // U+76E1 <cjk>
	0xE1B7: '盥' // U+76E5 <cjk>
	0xE1B8: '盧' // U+76E7 <cjk>
	0xE1B9: '盪' // U+76EA <cjk>
	0xE1BA: '蘯' // U+862F <cjk>
	0xE1BB: '盻' // U+76FB <cjk>
	0xE1BC: '眈' // U+7708 <cjk>
	0xE1BD: '眇' // U+7707 <cjk>
	0xE1BE: '眄' // U+7704 <cjk>
	0xE1BF: '眩' // U+7729 <cjk>
	0xE1C0: '眤' // U+7724 <cjk>
	0xE1C1: '眞' // U+771E <cjk>
	0xE1C2: '眥' // U+7725 <cjk>
	0xE1C3: '眦' // U+7726 <cjk>
	0xE1C4: '眛' // U+771B <cjk>
	0xE1C5: '眷' // U+7737 <cjk>
	0xE1C6: '眸' // U+7738 <cjk>
	0xE1C7: '睇' // U+7747 <cjk>
	0xE1C8: '睚' // U+775A <cjk>
	0xE1C9: '睨' // U+7768 <cjk>
	0xE1CA: '睫' // U+776B <cjk>
	0xE1CB: '睛' // U+775B <cjk>
	0xE1CC: '睥' // U+7765 <cjk>
	0xE1CD: '睿' // U+777F <cjk>
	0xE1CE: '睾' // U+777E <cjk>
	0xE1CF: '睹' // U+7779 <cjk>
	0xE1D0: '瞎' // U+778E <cjk>
	0xE1D1: '瞋' // U+778B <cjk>
	0xE1D2: '瞑' // U+7791 <cjk>
	0xE1D3: '瞠' // U+77A0 <cjk>
	0xE1D4: '瞞' // U+779E <cjk>
	0xE1D5: '瞰' // U+77B0 <cjk>
	0xE1D6: '瞶' // U+77B6 <cjk>
	0xE1D7: '瞹' // U+77B9 <cjk>
	0xE1D8: '瞿' // U+77BF <cjk>
	0xE1D9: '瞼' // U+77BC <cjk>
	0xE1DA: '瞽' // U+77BD <cjk>
	0xE1DB: '瞻' // U+77BB <cjk>
	0xE1DC: '矇' // U+77C7 <cjk>
	0xE1DD: '矍' // U+77CD <cjk>
	0xE1DE: '矗' // U+77D7 <cjk>
	0xE1DF: '矚' // U+77DA <cjk>
	0xE1E0: '矜' // U+77DC <cjk>
	0xE1E1: '矣' // U+77E3 <cjk>
	0xE1E2: '矮' // U+77EE <cjk>
	0xE1E3: '矼' // U+77FC <cjk>
	0xE1E4: '砌' // U+780C <cjk>
	0xE1E5: '砒' // U+7812 <cjk>
	0xE1E6: '礦' // U+7926 <cjk>
	0xE1E7: '砠' // U+7820 <cjk>
	0xE1E8: '礪' // U+792A <cjk>
	0xE1E9: '硅' // U+7845 <cjk>
	0xE1EA: '碎' // U+788E <cjk>
	0xE1EB: '硴' // U+7874 <cjk>
	0xE1EC: '碆' // U+7886 <cjk>
	0xE1ED: '硼' // U+787C <cjk>
	0xE1EE: '碚' // U+789A <cjk>
	0xE1EF: '碌' // U+788C <cjk>
	0xE1F0: '碣' // U+78A3 <cjk>
	0xE1F1: '碵' // U+78B5 <cjk>
	0xE1F2: '碪' // U+78AA <cjk>
	0xE1F3: '碯' // U+78AF <cjk>
	0xE1F4: '磑' // U+78D1 <cjk>
	0xE1F5: '磆' // U+78C6 <cjk>
	0xE1F6: '磋' // U+78CB <cjk>
	0xE1F7: '磔' // U+78D4 <cjk>
	0xE1F8: '碾' // U+78BE <cjk>
	0xE1F9: '碼' // U+78BC <cjk>
	0xE1FA: '磅' // U+78C5 <cjk>
	0xE1FB: '磊' // U+78CA <cjk>
	0xE1FC: '磬' // U+78EC <cjk>
	0xE240: '磧' // U+78E7 <cjk>
	0xE241: '磚' // U+78DA <cjk>
	0xE242: '磽' // U+78FD <cjk>
	0xE243: '磴' // U+78F4 <cjk>
	0xE244: '礇' // U+7907 <cjk>
	0xE245: '礒' // U+7912 <cjk>
	0xE246: '礑' // U+7911 <cjk>
	0xE247: '礙' // U+7919 <cjk>
	0xE248: '礬' // U+792C <cjk>
	0xE249: '礫' // U+792B <cjk>
	0xE24A: '祀' // U+7940 <cjk>
	0xE24B: '祠' // U+7960 <cjk>
	0xE24C: '祗' // U+7957 <cjk>
	0xE24D: '祟' // U+795F <cjk>
	0xE24E: '祚' // U+795A <cjk>
	0xE24F: '祕' // U+7955 <cjk>
	0xE250: '祓' // U+7953 <cjk>
	0xE251: '祺' // U+797A <cjk>
	0xE252: '祿' // U+797F <cjk>
	0xE253: '禊' // U+798A <cjk>
	0xE254: '禝' // U+799D <cjk>
	0xE255: '禧' // U+79A7 <cjk>
	0xE256: '齋' // U+9F4B <cjk>
	0xE257: '禪' // U+79AA <cjk>
	0xE258: '禮' // U+79AE <cjk>
	0xE259: '禳' // U+79B3 <cjk>
	0xE25A: '禹' // U+79B9 <cjk>
	0xE25B: '禺' // U+79BA <cjk>
	0xE25C: '秉' // U+79C9 <cjk>
	0xE25D: '秕' // U+79D5 <cjk>
	0xE25E: '秧' // U+79E7 <cjk>
	0xE25F: '秬' // U+79EC <cjk>
	0xE260: '秡' // U+79E1 <cjk>
	0xE261: '秣' // U+79E3 <cjk>
	0xE262: '稈' // U+7A08 <cjk>
	0xE263: '稍' // U+7A0D <cjk>
	0xE264: '稘' // U+7A18 <cjk>
	0xE265: '稙' // U+7A19 <cjk>
	0xE266: '稠' // U+7A20 <cjk>
	0xE267: '稟' // U+7A1F <cjk>
	0xE268: '禀' // U+7980 <cjk>
	0xE269: '稱' // U+7A31 <cjk>
	0xE26A: '稻' // U+7A3B <cjk>
	0xE26B: '稾' // U+7A3E <cjk>
	0xE26C: '稷' // U+7A37 <cjk>
	0xE26D: '穃' // U+7A43 <cjk>
	0xE26E: '穗' // U+7A57 <cjk>
	0xE26F: '穉' // U+7A49 <cjk>
	0xE270: '穡' // U+7A61 <cjk>
	0xE271: '穢' // U+7A62 <cjk>
	0xE272: '穩' // U+7A69 <cjk>
	0xE273: '龝' // U+9F9D <cjk>
	0xE274: '穰' // U+7A70 <cjk>
	0xE275: '穹' // U+7A79 <cjk>
	0xE276: '穽' // U+7A7D <cjk>
	0xE277: '窈' // U+7A88 <cjk>
	0xE278: '窗' // U+7A97 <cjk>
	0xE279: '窕' // U+7A95 <cjk>
	0xE27A: '窘' // U+7A98 <cjk>
	0xE27B: '窖' // U+7A96 <cjk>
	0xE27C: '窩' // U+7AA9 <cjk>
	0xE27D: '竈' // U+7AC8 <cjk>
	0xE27E: '窰' // U+7AB0 <cjk>
	0xE280: '窶' // U+7AB6 <cjk>
	0xE281: '竅' // U+7AC5 <cjk>
	0xE282: '竄' // U+7AC4 <cjk>
	0xE283: '窿' // U+7ABF <cjk>
	0xE284: '邃' // U+9083 <cjk>
	0xE285: '竇' // U+7AC7 <cjk>
	0xE286: '竊' // U+7ACA <cjk>
	0xE287: '竍' // U+7ACD <cjk>
	0xE288: '竏' // U+7ACF <cjk>
	0xE289: '竕' // U+7AD5 <cjk>
	0xE28A: '竓' // U+7AD3 <cjk>
	0xE28B: '站' // U+7AD9 <cjk>
	0xE28C: '竚' // U+7ADA <cjk>
	0xE28D: '竝' // U+7ADD <cjk>
	0xE28E: '竡' // U+7AE1 <cjk>
	0xE28F: '竢' // U+7AE2 <cjk>
	0xE290: '竦' // U+7AE6 <cjk>
	0xE291: '竭' // U+7AED <cjk>
	0xE292: '竰' // U+7AF0 <cjk>
	0xE293: '笂' // U+7B02 <cjk>
	0xE294: '笏' // U+7B0F <cjk>
	0xE295: '笊' // U+7B0A <cjk>
	0xE296: '笆' // U+7B06 <cjk>
	0xE297: '笳' // U+7B33 <cjk>
	0xE298: '笘' // U+7B18 <cjk>
	0xE299: '笙' // U+7B19 <cjk>
	0xE29A: '笞' // U+7B1E <cjk>
	0xE29B: '笵' // U+7B35 <cjk>
	0xE29C: '笨' // U+7B28 <cjk>
	0xE29D: '笶' // U+7B36 <cjk>
	0xE29E: '筐' // U+7B50 <cjk>
	0xE29F: '筺' // U+7B7A <cjk>
	0xE2A0: '笄' // U+7B04 <cjk>
	0xE2A1: '筍' // U+7B4D <cjk>
	0xE2A2: '笋' // U+7B0B <cjk>
	0xE2A3: '筌' // U+7B4C <cjk>
	0xE2A4: '筅' // U+7B45 <cjk>
	0xE2A5: '筵' // U+7B75 <cjk>
	0xE2A6: '筥' // U+7B65 <cjk>
	0xE2A7: '筴' // U+7B74 <cjk>
	0xE2A8: '筧' // U+7B67 <cjk>
	0xE2A9: '筰' // U+7B70 <cjk>
	0xE2AA: '筱' // U+7B71 <cjk>
	0xE2AB: '筬' // U+7B6C <cjk>
	0xE2AC: '筮' // U+7B6E <cjk>
	0xE2AD: '箝' // U+7B9D <cjk>
	0xE2AE: '箘' // U+7B98 <cjk>
	0xE2AF: '箟' // U+7B9F <cjk>
	0xE2B0: '箍' // U+7B8D <cjk>
	0xE2B1: '箜' // U+7B9C <cjk>
	0xE2B2: '箚' // U+7B9A <cjk>
	0xE2B3: '箋' // U+7B8B <cjk>
	0xE2B4: '箒' // U+7B92 <cjk>
	0xE2B5: '箏' // U+7B8F <cjk>
	0xE2B6: '筝' // U+7B5D <cjk>
	0xE2B7: '箙' // U+7B99 <cjk>
	0xE2B8: '篋' // U+7BCB <cjk>
	0xE2B9: '篁' // U+7BC1 <cjk>
	0xE2BA: '篌' // U+7BCC <cjk>
	0xE2BB: '篏' // U+7BCF <cjk>
	0xE2BC: '箴' // U+7BB4 <cjk>
	0xE2BD: '篆' // U+7BC6 <cjk>
	0xE2BE: '篝' // U+7BDD <cjk>
	0xE2BF: '篩' // U+7BE9 <cjk>
	0xE2C0: '簑' // U+7C11 <cjk>
	0xE2C1: '簔' // U+7C14 <cjk>
	0xE2C2: '篦' // U+7BE6 <cjk>
	0xE2C3: '篥' // U+7BE5 <cjk>
	0xE2C4: '籠' // U+7C60 <cjk>
	0xE2C5: '簀' // U+7C00 <cjk>
	0xE2C6: '簇' // U+7C07 <cjk>
	0xE2C7: '簓' // U+7C13 <cjk>
	0xE2C8: '篳' // U+7BF3 <cjk>
	0xE2C9: '篷' // U+7BF7 <cjk>
	0xE2CA: '簗' // U+7C17 <cjk>
	0xE2CB: '簍' // U+7C0D <cjk>
	0xE2CC: '篶' // U+7BF6 <cjk>
	0xE2CD: '簣' // U+7C23 <cjk>
	0xE2CE: '簧' // U+7C27 <cjk>
	0xE2CF: '簪' // U+7C2A <cjk>
	0xE2D0: '簟' // U+7C1F <cjk>
	0xE2D1: '簷' // U+7C37 <cjk>
	0xE2D2: '簫' // U+7C2B <cjk>
	0xE2D3: '簽' // U+7C3D <cjk>
	0xE2D4: '籌' // U+7C4C <cjk>
	0xE2D5: '籃' // U+7C43 <cjk>
	0xE2D6: '籔' // U+7C54 <cjk>
	0xE2D7: '籏' // U+7C4F <cjk>
	0xE2D8: '籀' // U+7C40 <cjk>
	0xE2D9: '籐' // U+7C50 <cjk>
	0xE2DA: '籘' // U+7C58 <cjk>
	0xE2DB: '籟' // U+7C5F <cjk>
	0xE2DC: '籤' // U+7C64 <cjk>
	0xE2DD: '籖' // U+7C56 <cjk>
	0xE2DE: '籥' // U+7C65 <cjk>
	0xE2DF: '籬' // U+7C6C <cjk>
	0xE2E0: '籵' // U+7C75 <cjk>
	0xE2E1: '粃' // U+7C83 <cjk>
	0xE2E2: '粐' // U+7C90 <cjk>
	0xE2E3: '粤' // U+7CA4 <cjk>
	0xE2E4: '粭' // U+7CAD <cjk>
	0xE2E5: '粢' // U+7CA2 <cjk>
	0xE2E6: '粫' // U+7CAB <cjk>
	0xE2E7: '粡' // U+7CA1 <cjk>
	0xE2E8: '粨' // U+7CA8 <cjk>
	0xE2E9: '粳' // U+7CB3 <cjk>
	0xE2EA: '粲' // U+7CB2 <cjk>
	0xE2EB: '粱' // U+7CB1 <cjk>
	0xE2EC: '粮' // U+7CAE <cjk>
	0xE2ED: '粹' // U+7CB9 <cjk>
	0xE2EE: '粽' // U+7CBD <cjk>
	0xE2EF: '糀' // U+7CC0 <cjk>
	0xE2F0: '糅' // U+7CC5 <cjk>
	0xE2F1: '糂' // U+7CC2 <cjk>
	0xE2F2: '糘' // U+7CD8 <cjk>
	0xE2F3: '糒' // U+7CD2 <cjk>
	0xE2F4: '糜' // U+7CDC <cjk>
	0xE2F5: '糢' // U+7CE2 <cjk>
	0xE2F6: '鬻' // U+9B3B <cjk>
	0xE2F7: '糯' // U+7CEF <cjk>
	0xE2F8: '糲' // U+7CF2 <cjk>
	0xE2F9: '糴' // U+7CF4 <cjk>
	0xE2FA: '糶' // U+7CF6 <cjk>
	0xE2FB: '糺' // U+7CFA <cjk>
	0xE2FC: '紆' // U+7D06 <cjk>
	0xE340: '紂' // U+7D02 <cjk>
	0xE341: '紜' // U+7D1C <cjk>
	0xE342: '紕' // U+7D15 <cjk>
	0xE343: '紊' // U+7D0A <cjk>
	0xE344: '絅' // U+7D45 <cjk>
	0xE345: '絋' // U+7D4B <cjk>
	0xE346: '紮' // U+7D2E <cjk>
	0xE347: '紲' // U+7D32 <cjk>
	0xE348: '紿' // U+7D3F <cjk>
	0xE349: '紵' // U+7D35 <cjk>
	0xE34A: '絆' // U+7D46 <cjk>
	0xE34B: '絳' // U+7D73 <cjk>
	0xE34C: '絖' // U+7D56 <cjk>
	0xE34D: '絎' // U+7D4E <cjk>
	0xE34E: '絲' // U+7D72 <cjk>
	0xE34F: '絨' // U+7D68 <cjk>
	0xE350: '絮' // U+7D6E <cjk>
	0xE351: '絏' // U+7D4F <cjk>
	0xE352: '絣' // U+7D63 <cjk>
	0xE353: '經' // U+7D93 <cjk>
	0xE354: '綉' // U+7D89 <cjk>
	0xE355: '絛' // U+7D5B <cjk>
	0xE356: '綏' // U+7D8F <cjk>
	0xE357: '絽' // U+7D7D <cjk>
	0xE358: '綛' // U+7D9B <cjk>
	0xE359: '綺' // U+7DBA <cjk>
	0xE35A: '綮' // U+7DAE <cjk>
	0xE35B: '綣' // U+7DA3 <cjk>
	0xE35C: '綵' // U+7DB5 <cjk>
	0xE35D: '緇' // U+7DC7 <cjk>
	0xE35E: '綽' // U+7DBD <cjk>
	0xE35F: '綫' // U+7DAB <cjk>
	0xE360: '總' // U+7E3D <cjk>
	0xE361: '綢' // U+7DA2 <cjk>
	0xE362: '綯' // U+7DAF <cjk>
	0xE363: '緜' // U+7DDC <cjk>
	0xE364: '綸' // U+7DB8 <cjk>
	0xE365: '綟' // U+7D9F <cjk>
	0xE366: '綰' // U+7DB0 <cjk>
	0xE367: '緘' // U+7DD8 <cjk>
	0xE368: '緝' // U+7DDD <cjk>
	0xE369: '緤' // U+7DE4 <cjk>
	0xE36A: '緞' // U+7DDE <cjk>
	0xE36B: '緻' // U+7DFB <cjk>
	0xE36C: '緲' // U+7DF2 <cjk>
	0xE36D: '緡' // U+7DE1 <cjk>
	0xE36E: '縅' // U+7E05 <cjk>
	0xE36F: '縊' // U+7E0A <cjk>
	0xE370: '縣' // U+7E23 <cjk>
	0xE371: '縡' // U+7E21 <cjk>
	0xE372: '縒' // U+7E12 <cjk>
	0xE373: '縱' // U+7E31 <cjk>
	0xE374: '縟' // U+7E1F <cjk>
	0xE375: '縉' // U+7E09 <cjk>
	0xE376: '縋' // U+7E0B <cjk>
	0xE377: '縢' // U+7E22 <cjk>
	0xE378: '繆' // U+7E46 <cjk>
	0xE379: '繦' // U+7E66 <cjk>
	0xE37A: '縻' // U+7E3B <cjk>
	0xE37B: '縵' // U+7E35 <cjk>
	0xE37C: '縹' // U+7E39 <cjk>
	0xE37D: '繃' // U+7E43 <cjk>
	0xE37E: '縷' // U+7E37 <cjk>
	0xE380: '縲' // U+7E32 <cjk>
	0xE381: '縺' // U+7E3A <cjk>
	0xE382: '繧' // U+7E67 <cjk>
	0xE383: '繝' // U+7E5D <cjk>
	0xE384: '繖' // U+7E56 <cjk>
	0xE385: '繞' // U+7E5E <cjk>
	0xE386: '繙' // U+7E59 <cjk>
	0xE387: '繚' // U+7E5A <cjk>
	0xE388: '繹' // U+7E79 <cjk>
	0xE389: '繪' // U+7E6A <cjk>
	0xE38A: '繩' // U+7E69 <cjk>
	0xE38B: '繼' // U+7E7C <cjk>
	0xE38C: '繻' // U+7E7B <cjk>
	0xE38D: '纃' // U+7E83 <cjk>
	0xE38E: '緕' // U+7DD5 <cjk>
	0xE38F: '繽' // U+7E7D <cjk>
	0xE390: '辮' // U+8FAE <cjk>
	0xE391: '繿' // U+7E7F <cjk>
	0xE392: '纈' // U+7E88 <cjk>
	0xE393: '纉' // U+7E89 <cjk>
	0xE394: '續' // U+7E8C <cjk>
	0xE395: '纒' // U+7E92 <cjk>
	0xE396: '纐' // U+7E90 <cjk>
	0xE397: '纓' // U+7E93 <cjk>
	0xE398: '纔' // U+7E94 <cjk>
	0xE399: '纖' // U+7E96 <cjk>
	0xE39A: '纎' // U+7E8E <cjk>
	0xE39B: '纛' // U+7E9B <cjk>
	0xE39C: '纜' // U+7E9C <cjk>
	0xE39D: '缸' // U+7F38 <cjk>
	0xE39E: '缺' // U+7F3A <cjk>
	0xE39F: '罅' // U+7F45 <cjk>
	0xE3A0: '罌' // U+7F4C <cjk>
	0xE3A1: '罍' // U+7F4D <cjk>
	0xE3A2: '罎' // U+7F4E <cjk>
	0xE3A3: '罐' // U+7F50 <cjk>
	0xE3A4: '网' // U+7F51 <cjk>
	0xE3A5: '罕' // U+7F55 <cjk>
	0xE3A6: '罔' // U+7F54 <cjk>
	0xE3A7: '罘' // U+7F58 <cjk>
	0xE3A8: '罟' // U+7F5F <cjk>
	0xE3A9: '罠' // U+7F60 <cjk>
	0xE3AA: '罨' // U+7F68 <cjk>
	0xE3AB: '罩' // U+7F69 <cjk>
	0xE3AC: '罧' // U+7F67 <cjk>
	0xE3AD: '罸' // U+7F78 <cjk>
	0xE3AE: '羂' // U+7F82 <cjk>
	0xE3AF: '羆' // U+7F86 <cjk>
	0xE3B0: '羃' // U+7F83 <cjk>
	0xE3B1: '羈' // U+7F88 <cjk>
	0xE3B2: '羇' // U+7F87 <cjk>
	0xE3B3: '羌' // U+7F8C <cjk>
	0xE3B4: '羔' // U+7F94 <cjk>
	0xE3B5: '羞' // U+7F9E <cjk>
	0xE3B6: '羝' // U+7F9D <cjk>
	0xE3B7: '羚' // U+7F9A <cjk>
	0xE3B8: '羣' // U+7FA3 <cjk>
	0xE3B9: '羯' // U+7FAF <cjk>
	0xE3BA: '羲' // U+7FB2 <cjk>
	0xE3BB: '羹' // U+7FB9 <cjk>
	0xE3BC: '羮' // U+7FAE <cjk>
	0xE3BD: '羶' // U+7FB6 <cjk>
	0xE3BE: '羸' // U+7FB8 <cjk>
	0xE3BF: '譱' // U+8B71 <cjk>
	0xE3C0: '翅' // U+7FC5 <cjk>
	0xE3C1: '翆' // U+7FC6 <cjk>
	0xE3C2: '翊' // U+7FCA <cjk>
	0xE3C3: '翕' // U+7FD5 <cjk>
	0xE3C4: '翔' // U+7FD4 <cjk>
	0xE3C5: '翡' // U+7FE1 <cjk>
	0xE3C6: '翦' // U+7FE6 <cjk>
	0xE3C7: '翩' // U+7FE9 <cjk>
	0xE3C8: '翳' // U+7FF3 <cjk>
	0xE3C9: '翹' // U+7FF9 <cjk>
	0xE3CA: '飜' // U+98DC <cjk>
	0xE3CB: '耆' // U+8006 <cjk>
	0xE3CC: '耄' // U+8004 <cjk>
	0xE3CD: '耋' // U+800B <cjk>
	0xE3CE: '耒' // U+8012 <cjk>
	0xE3CF: '耘' // U+8018 <cjk>
	0xE3D0: '耙' // U+8019 <cjk>
	0xE3D1: '耜' // U+801C <cjk>
	0xE3D2: '耡' // U+8021 <cjk>
	0xE3D3: '耨' // U+8028 <cjk>
	0xE3D4: '耿' // U+803F <cjk>
	0xE3D5: '耻' // U+803B <cjk>
	0xE3D6: '聊' // U+804A <cjk>
	0xE3D7: '聆' // U+8046 <cjk>
	0xE3D8: '聒' // U+8052 <cjk>
	0xE3D9: '聘' // U+8058 <cjk>
	0xE3DA: '聚' // U+805A <cjk>
	0xE3DB: '聟' // U+805F <cjk>
	0xE3DC: '聢' // U+8062 <cjk>
	0xE3DD: '聨' // U+8068 <cjk>
	0xE3DE: '聳' // U+8073 <cjk>
	0xE3DF: '聲' // U+8072 <cjk>
	0xE3E0: '聰' // U+8070 <cjk>
	0xE3E1: '聶' // U+8076 <cjk>
	0xE3E2: '聹' // U+8079 <cjk>
	0xE3E3: '聽' // U+807D <cjk>
	0xE3E4: '聿' // U+807F <cjk>
	0xE3E5: '肄' // U+8084 <cjk>
	0xE3E6: '肆' // U+8086 <cjk>
	0xE3E7: '肅' // U+8085 <cjk>
	0xE3E8: '肛' // U+809B <cjk>
	0xE3E9: '肓' // U+8093 <cjk>
	0xE3EA: '肚' // U+809A <cjk>
	0xE3EB: '肭' // U+80AD <cjk>
	0xE3EC: '冐' // U+5190 <cjk>
	0xE3ED: '肬' // U+80AC <cjk>
	0xE3EE: '胛' // U+80DB <cjk>
	0xE3EF: '胥' // U+80E5 <cjk>
	0xE3F0: '胙' // U+80D9 <cjk>
	0xE3F1: '胝' // U+80DD <cjk>
	0xE3F2: '胄' // U+80C4 <cjk>
	0xE3F3: '胚' // U+80DA <cjk>
	0xE3F4: '胖' // U+80D6 <cjk>
	0xE3F5: '脉' // U+8109 <cjk>
	0xE3F6: '胯' // U+80EF <cjk>
	0xE3F7: '胱' // U+80F1 <cjk>
	0xE3F8: '脛' // U+811B <cjk>
	0xE3F9: '脩' // U+8129 <cjk>
	0xE3FA: '脣' // U+8123 <cjk>
	0xE3FB: '脯' // U+812F <cjk>
	0xE3FC: '腋' // U+814B <cjk>
	0xE440: '隋' // U+968B <cjk>
	0xE441: '腆' // U+8146 <cjk>
	0xE442: '脾' // U+813E <cjk>
	0xE443: '腓' // U+8153 <cjk>
	0xE444: '腑' // U+8151 <cjk>
	0xE445: '胼' // U+80FC <cjk>
	0xE446: '腱' // U+8171 <cjk>
	0xE447: '腮' // U+816E <cjk>
	0xE448: '腥' // U+8165 <cjk>
	0xE449: '腦' // U+8166 <cjk>
	0xE44A: '腴' // U+8174 <cjk>
	0xE44B: '膃' // U+8183 <cjk>
	0xE44C: '膈' // U+8188 <cjk>
	0xE44D: '膊' // U+818A <cjk>
	0xE44E: '膀' // U+8180 <cjk>
	0xE44F: '膂' // U+8182 <cjk>
	0xE450: '膠' // U+81A0 <cjk>
	0xE451: '膕' // U+8195 <cjk>
	0xE452: '膤' // U+81A4 <cjk>
	0xE453: '膣' // U+81A3 <cjk>
	0xE454: '腟' // U+815F <cjk>
	0xE455: '膓' // U+8193 <cjk>
	0xE456: '膩' // U+81A9 <cjk>
	0xE457: '膰' // U+81B0 <cjk>
	0xE458: '膵' // U+81B5 <cjk>
	0xE459: '膾' // U+81BE <cjk>
	0xE45A: '膸' // U+81B8 <cjk>
	0xE45B: '膽' // U+81BD <cjk>
	0xE45C: '臀' // U+81C0 <cjk>
	0xE45D: '臂' // U+81C2 <cjk>
	0xE45E: '膺' // U+81BA <cjk>
	0xE45F: '臉' // U+81C9 <cjk>
	0xE460: '臍' // U+81CD <cjk>
	0xE461: '臑' // U+81D1 <cjk>
	0xE462: '臙' // U+81D9 <cjk>
	0xE463: '臘' // U+81D8 <cjk>
	0xE464: '臈' // U+81C8 <cjk>
	0xE465: '臚' // U+81DA <cjk>
	0xE466: '臟' // U+81DF <cjk>
	0xE467: '臠' // U+81E0 <cjk>
	0xE468: '臧' // U+81E7 <cjk>
	0xE469: '臺' // U+81FA <cjk>
	0xE46A: '臻' // U+81FB <cjk>
	0xE46B: '臾' // U+81FE <cjk>
	0xE46C: '舁' // U+8201 <cjk>
	0xE46D: '舂' // U+8202 <cjk>
	0xE46E: '舅' // U+8205 <cjk>
	0xE46F: '與' // U+8207 <cjk>
	0xE470: '舊' // U+820A <cjk>
	0xE471: '舍' // U+820D <cjk>
	0xE472: '舐' // U+8210 <cjk>
	0xE473: '舖' // U+8216 <cjk>
	0xE474: '舩' // U+8229 <cjk>
	0xE475: '舫' // U+822B <cjk>
	0xE476: '舸' // U+8238 <cjk>
	0xE477: '舳' // U+8233 <cjk>
	0xE478: '艀' // U+8240 <cjk>
	0xE479: '艙' // U+8259 <cjk>
	0xE47A: '艘' // U+8258 <cjk>
	0xE47B: '艝' // U+825D <cjk>
	0xE47C: '艚' // U+825A <cjk>
	0xE47D: '艟' // U+825F <cjk>
	0xE47E: '艤' // U+8264 <cjk>
	0xE480: '艢' // U+8262 <cjk>
	0xE481: '艨' // U+8268 <cjk>
	0xE482: '艪' // U+826A <cjk>
	0xE483: '艫' // U+826B <cjk>
	0xE484: '舮' // U+822E <cjk>
	0xE485: '艱' // U+8271 <cjk>
	0xE486: '艷' // U+8277 <cjk>
	0xE487: '艸' // U+8278 <cjk>
	0xE488: '艾' // U+827E <cjk>
	0xE489: '芍' // U+828D <cjk>
	0xE48A: '芒' // U+8292 <cjk>
	0xE48B: '芫' // U+82AB <cjk>
	0xE48C: '芟' // U+829F <cjk>
	0xE48D: '芻' // U+82BB <cjk>
	0xE48E: '芬' // U+82AC <cjk>
	0xE48F: '苡' // U+82E1 <cjk>
	0xE490: '苣' // U+82E3 <cjk>
	0xE491: '苟' // U+82DF <cjk>
	0xE492: '苒' // U+82D2 <cjk>
	0xE493: '苴' // U+82F4 <cjk>
	0xE494: '苳' // U+82F3 <cjk>
	0xE495: '苺' // U+82FA <cjk>
	0xE496: '莓' // U+8393 <cjk>
	0xE497: '范' // U+8303 <cjk>
	0xE498: '苻' // U+82FB <cjk>
	0xE499: '苹' // U+82F9 <cjk>
	0xE49A: '苞' // U+82DE <cjk>
	0xE49B: '茆' // U+8306 <cjk>
	0xE49C: '苜' // U+82DC <cjk>
	0xE49D: '茉' // U+8309 <cjk>
	0xE49E: '苙' // U+82D9 <cjk>
	0xE49F: '茵' // U+8335 <cjk>
	0xE4A0: '茴' // U+8334 <cjk>
	0xE4A1: '茖' // U+8316 <cjk>
	0xE4A2: '茲' // U+8332 <cjk>
	0xE4A3: '茱' // U+8331 <cjk>
	0xE4A4: '荀' // U+8340 <cjk>
	0xE4A5: '茹' // U+8339 <cjk>
	0xE4A6: '荐' // U+8350 <cjk>
	0xE4A7: '荅' // U+8345 <cjk>
	0xE4A8: '茯' // U+832F <cjk>
	0xE4A9: '茫' // U+832B <cjk>
	0xE4AA: '茗' // U+8317 <cjk>
	0xE4AB: '茘' // U+8318 <cjk>
	0xE4AC: '莅' // U+8385 <cjk>
	0xE4AD: '莚' // U+839A <cjk>
	0xE4AE: '莪' // U+83AA <cjk>
	0xE4AF: '莟' // U+839F <cjk>
	0xE4B0: '莢' // U+83A2 <cjk>
	0xE4B1: '莖' // U+8396 <cjk>
	0xE4B2: '茣' // U+8323 <cjk>
	0xE4B3: '莎' // U+838E <cjk>
	0xE4B4: '莇' // U+8387 <cjk>
	0xE4B5: '莊' // U+838A <cjk>
	0xE4B6: '荼' // U+837C <cjk>
	0xE4B7: '莵' // U+83B5 <cjk>
	0xE4B8: '荳' // U+8373 <cjk>
	0xE4B9: '荵' // U+8375 <cjk>
	0xE4BA: '莠' // U+83A0 <cjk>
	0xE4BB: '莉' // U+8389 <cjk>
	0xE4BC: '莨' // U+83A8 <cjk>
	0xE4BD: '菴' // U+83F4 <cjk>
	0xE4BE: '萓' // U+8413 <cjk>
	0xE4BF: '菫' // U+83EB <cjk>
	0xE4C0: '菎' // U+83CE <cjk>
	0xE4C1: '菽' // U+83FD <cjk>
	0xE4C2: '萃' // U+8403 <cjk>
	0xE4C3: '菘' // U+83D8 <cjk>
	0xE4C4: '萋' // U+840B <cjk>
	0xE4C5: '菁' // U+83C1 <cjk>
	0xE4C6: '菷' // U+83F7 <cjk>
	0xE4C7: '萇' // U+8407 <cjk>
	0xE4C8: '菠' // U+83E0 <cjk>
	0xE4C9: '菲' // U+83F2 <cjk>
	0xE4CA: '萍' // U+840D <cjk>
	0xE4CB: '萢' // U+8422 <cjk>
	0xE4CC: '萠' // U+8420 <cjk>
	0xE4CD: '莽' // U+83BD <cjk>
	0xE4CE: '萸' // U+8438 <cjk>
	0xE4CF: '蔆' // U+8506 <cjk>
	0xE4D0: '菻' // U+83FB <cjk>
	0xE4D1: '葭' // U+846D <cjk>
	0xE4D2: '萪' // U+842A <cjk>
	0xE4D3: '萼' // U+843C <cjk>
	0xE4D4: '蕚' // U+855A <cjk>
	0xE4D5: '蒄' // U+8484 <cjk>
	0xE4D6: '葷' // U+8477 <cjk>
	0xE4D7: '葫' // U+846B <cjk>
	0xE4D8: '蒭' // U+84AD <cjk>
	0xE4D9: '葮' // U+846E <cjk>
	0xE4DA: '蒂' // U+8482 <cjk>
	0xE4DB: '葩' // U+8469 <cjk>
	0xE4DC: '葆' // U+8446 <cjk>
	0xE4DD: '萬' // U+842C <cjk>
	0xE4DE: '葯' // U+846F <cjk>
	0xE4DF: '葹' // U+8479 <cjk>
	0xE4E0: '萵' // U+8435 <cjk>
	0xE4E1: '蓊' // U+84CA <cjk>
	0xE4E2: '葢' // U+8462 <cjk>
	0xE4E3: '蒹' // U+84B9 <cjk>
	0xE4E4: '蒿' // U+84BF <cjk>
	0xE4E5: '蒟' // U+849F <cjk>
	0xE4E6: '蓙' // U+84D9 <cjk>
	0xE4E7: '蓍' // U+84CD <cjk>
	0xE4E8: '蒻' // U+84BB <cjk>
	0xE4E9: '蓚' // U+84DA <cjk>
	0xE4EA: '蓐' // U+84D0 <cjk>
	0xE4EB: '蓁' // U+84C1 <cjk>
	0xE4EC: '蓆' // U+84C6 <cjk>
	0xE4ED: '蓖' // U+84D6 <cjk>
	0xE4EE: '蒡' // U+84A1 <cjk>
	0xE4EF: '蔡' // U+8521 <cjk>
	0xE4F0: '蓿' // U+84FF <cjk>
	0xE4F1: '蓴' // U+84F4 <cjk>
	0xE4F2: '蔗' // U+8517 <cjk>
	0xE4F3: '蔘' // U+8518 <cjk>
	0xE4F4: '蔬' // U+852C <cjk>
	0xE4F5: '蔟' // U+851F <cjk>
	0xE4F6: '蔕' // U+8515 <cjk>
	0xE4F7: '蔔' // U+8514 <cjk>
	0xE4F8: '蓼' // U+84FC <cjk>
	0xE4F9: '蕀' // U+8540 <cjk>
	0xE4FA: '蕣' // U+8563 <cjk>
	0xE4FB: '蕘' // U+8558 <cjk>
	0xE4FC: '蕈' // U+8548 <cjk>
	0xE540: '蕁' // U+8541 <cjk>
	0xE541: '蘂' // U+8602 <cjk>
	0xE542: '蕋' // U+854B <cjk>
	0xE543: '蕕' // U+8555 <cjk>
	0xE544: '薀' // U+8580 <cjk>
	0xE545: '薤' // U+85A4 <cjk>
	0xE546: '薈' // U+8588 <cjk>
	0xE547: '薑' // U+8591 <cjk>
	0xE548: '薊' // U+858A <cjk>
	0xE549: '薨' // U+85A8 <cjk>
	0xE54A: '蕭' // U+856D <cjk>
	0xE54B: '薔' // U+8594 <cjk>
	0xE54C: '薛' // U+859B <cjk>
	0xE54D: '藪' // U+85EA <cjk>
	0xE54E: '薇' // U+8587 <cjk>
	0xE54F: '薜' // U+859C <cjk>
	0xE550: '蕷' // U+8577 <cjk>
	0xE551: '蕾' // U+857E <cjk>
	0xE552: '薐' // U+8590 <cjk>
	0xE553: '藉' // U+85C9 <cjk>
	0xE554: '薺' // U+85BA <cjk>
	0xE555: '藏' // U+85CF <cjk>
	0xE556: '薹' // U+85B9 <cjk>
	0xE557: '藐' // U+85D0 <cjk>
	0xE558: '藕' // U+85D5 <cjk>
	0xE559: '藝' // U+85DD <cjk>
	0xE55A: '藥' // U+85E5 <cjk>
	0xE55B: '藜' // U+85DC <cjk>
	0xE55C: '藹' // U+85F9 <cjk>
	0xE55D: '蘊' // U+860A <cjk>
	0xE55E: '蘓' // U+8613 <cjk>
	0xE55F: '蘋' // U+860B <cjk>
	0xE560: '藾' // U+85FE <cjk>
	0xE561: '藺' // U+85FA <cjk>
	0xE562: '蘆' // U+8606 <cjk>
	0xE563: '蘢' // U+8622 <cjk>
	0xE564: '蘚' // U+861A <cjk>
	0xE565: '蘰' // U+8630 <cjk>
	0xE566: '蘿' // U+863F <cjk>
	0xE567: '虍' // U+864D <cjk>
	0xE568: '乕' // U+4E55 <cjk>
	0xE569: '虔' // U+8654 <cjk>
	0xE56A: '號' // U+865F <cjk>
	0xE56B: '虧' // U+8667 <cjk>
	0xE56C: '虱' // U+8671 <cjk>
	0xE56D: '蚓' // U+8693 <cjk>
	0xE56E: '蚣' // U+86A3 <cjk>
	0xE56F: '蚩' // U+86A9 <cjk>
	0xE570: '蚪' // U+86AA <cjk>
	0xE571: '蚋' // U+868B <cjk>
	0xE572: '蚌' // U+868C <cjk>
	0xE573: '蚶' // U+86B6 <cjk>
	0xE574: '蚯' // U+86AF <cjk>
	0xE575: '蛄' // U+86C4 <cjk>
	0xE576: '蛆' // U+86C6 <cjk>
	0xE577: '蚰' // U+86B0 <cjk>
	0xE578: '蛉' // U+86C9 <cjk>
	0xE579: '蠣' // U+8823 <cjk>
	0xE57A: '蚫' // U+86AB <cjk>
	0xE57B: '蛔' // U+86D4 <cjk>
	0xE57C: '蛞' // U+86DE <cjk>
	0xE57D: '蛩' // U+86E9 <cjk>
	0xE57E: '蛬' // U+86EC <cjk>
	0xE580: '蛟' // U+86DF <cjk>
	0xE581: '蛛' // U+86DB <cjk>
	0xE582: '蛯' // U+86EF <cjk>
	0xE583: '蜒' // U+8712 <cjk>
	0xE584: '蜆' // U+8706 <cjk>
	0xE585: '蜈' // U+8708 <cjk>
	0xE586: '蜀' // U+8700 <cjk>
	0xE587: '蜃' // U+8703 <cjk>
	0xE588: '蛻' // U+86FB <cjk>
	0xE589: '蜑' // U+8711 <cjk>
	0xE58A: '蜉' // U+8709 <cjk>
	0xE58B: '蜍' // U+870D <cjk>
	0xE58C: '蛹' // U+86F9 <cjk>
	0xE58D: '蜊' // U+870A <cjk>
	0xE58E: '蜴' // U+8734 <cjk>
	0xE58F: '蜿' // U+873F <cjk>
	0xE590: '蜷' // U+8737 <cjk>
	0xE591: '蜻' // U+873B <cjk>
	0xE592: '蜥' // U+8725 <cjk>
	0xE593: '蜩' // U+8729 <cjk>
	0xE594: '蜚' // U+871A <cjk>
	0xE595: '蝠' // U+8760 <cjk>
	0xE596: '蝟' // U+875F <cjk>
	0xE597: '蝸' // U+8778 <cjk>
	0xE598: '蝌' // U+874C <cjk>
	0xE599: '蝎' // U+874E <cjk>
	0xE59A: '蝴' // U+8774 <cjk>
	0xE59B: '蝗' // U+8757 <cjk>
	0xE59C: '蝨' // U+8768 <cjk>
	0xE59D: '蝮' // U+876E <cjk>
	0xE59E: '蝙' // U+8759 <cjk>
	0xE59F: '蝓' // U+8753 <cjk>
	0xE5A0: '蝣' // U+8763 <cjk>
	0xE5A1: '蝪' // U+876A <cjk>
	0xE5A2: '蠅' // U+8805 <cjk>
	0xE5A3: '螢' // U+87A2 <cjk>
	0xE5A4: '螟' // U+879F <cjk>
	0xE5A5: '螂' // U+8782 <cjk>
	0xE5A6: '螯' // U+87AF <cjk>
	0xE5A7: '蟋' // U+87CB <cjk>
	0xE5A8: '螽' // U+87BD <cjk>
	0xE5A9: '蟀' // U+87C0 <cjk>
	0xE5AA: '蟐' // U+87D0 <cjk>
	0xE5AB: '雖' // U+96D6 <cjk>
	0xE5AC: '螫' // U+87AB <cjk>
	0xE5AD: '蟄' // U+87C4 <cjk>
	0xE5AE: '螳' // U+87B3 <cjk>
	0xE5AF: '蟇' // U+87C7 <cjk>
	0xE5B0: '蟆' // U+87C6 <cjk>
	0xE5B1: '螻' // U+87BB <cjk>
	0xE5B2: '蟯' // U+87EF <cjk>
	0xE5B3: '蟲' // U+87F2 <cjk>
	0xE5B4: '蟠' // U+87E0 <cjk>
	0xE5B5: '蠏' // U+880F <cjk>
	0xE5B6: '蠍' // U+880D <cjk>
	0xE5B7: '蟾' // U+87FE <cjk>
	0xE5B8: '蟶' // U+87F6 <cjk>
	0xE5B9: '蟷' // U+87F7 <cjk>
	0xE5BA: '蠎' // U+880E <cjk>
	0xE5BB: '蟒' // U+87D2 <cjk>
	0xE5BC: '蠑' // U+8811 <cjk>
	0xE5BD: '蠖' // U+8816 <cjk>
	0xE5BE: '蠕' // U+8815 <cjk>
	0xE5BF: '蠢' // U+8822 <cjk>
	0xE5C0: '蠡' // U+8821 <cjk>
	0xE5C1: '蠱' // U+8831 <cjk>
	0xE5C2: '蠶' // U+8836 <cjk>
	0xE5C3: '蠹' // U+8839 <cjk>
	0xE5C4: '蠧' // U+8827 <cjk>
	0xE5C5: '蠻' // U+883B <cjk>
	0xE5C6: '衄' // U+8844 <cjk>
	0xE5C7: '衂' // U+8842 <cjk>
	0xE5C8: '衒' // U+8852 <cjk>
	0xE5C9: '衙' // U+8859 <cjk>
	0xE5CA: '衞' // U+885E <cjk>
	0xE5CB: '衢' // U+8862 <cjk>
	0xE5CC: '衫' // U+886B <cjk>
	0xE5CD: '袁' // U+8881 <cjk>
	0xE5CE: '衾' // U+887E <cjk>
	0xE5CF: '袞' // U+889E <cjk>
	0xE5D0: '衵' // U+8875 <cjk>
	0xE5D1: '衽' // U+887D <cjk>
	0xE5D2: '袵' // U+88B5 <cjk>
	0xE5D3: '衲' // U+8872 <cjk>
	0xE5D4: '袂' // U+8882 <cjk>
	0xE5D5: '袗' // U+8897 <cjk>
	0xE5D6: '袒' // U+8892 <cjk>
	0xE5D7: '袮' // U+88AE <cjk>
	0xE5D8: '袙' // U+8899 <cjk>
	0xE5D9: '袢' // U+88A2 <cjk>
	0xE5DA: '袍' // U+888D <cjk>
	0xE5DB: '袤' // U+88A4 <cjk>
	0xE5DC: '袰' // U+88B0 <cjk>
	0xE5DD: '袿' // U+88BF <cjk>
	0xE5DE: '袱' // U+88B1 <cjk>
	0xE5DF: '裃' // U+88C3 <cjk>
	0xE5E0: '裄' // U+88C4 <cjk>
	0xE5E1: '裔' // U+88D4 <cjk>
	0xE5E2: '裘' // U+88D8 <cjk>
	0xE5E3: '裙' // U+88D9 <cjk>
	0xE5E4: '裝' // U+88DD <cjk>
	0xE5E5: '裹' // U+88F9 <cjk>
	0xE5E6: '褂' // U+8902 <cjk>
	0xE5E7: '裼' // U+88FC <cjk>
	0xE5E8: '裴' // U+88F4 <cjk>
	0xE5E9: '裨' // U+88E8 <cjk>
	0xE5EA: '裲' // U+88F2 <cjk>
	0xE5EB: '褄' // U+8904 <cjk>
	0xE5EC: '褌' // U+890C <cjk>
	0xE5ED: '褊' // U+890A <cjk>
	0xE5EE: '褓' // U+8913 <cjk>
	0xE5EF: '襃' // U+8943 <cjk>
	0xE5F0: '褞' // U+891E <cjk>
	0xE5F1: '褥' // U+8925 <cjk>
	0xE5F2: '褪' // U+892A <cjk>
	0xE5F3: '褫' // U+892B <cjk>
	0xE5F4: '襁' // U+8941 <cjk>
	0xE5F5: '襄' // U+8944 <cjk>
	0xE5F6: '褻' // U+893B <cjk>
	0xE5F7: '褶' // U+8936 <cjk>
	0xE5F8: '褸' // U+8938 <cjk>
	0xE5F9: '襌' // U+894C <cjk>
	0xE5FA: '褝' // U+891D <cjk>
	0xE5FB: '襠' // U+8960 <cjk>
	0xE5FC: '襞' // U+895E <cjk>
	0xE640: '襦' // U+8966 <cjk>
	0xE641: '襤' // U+8964 <cjk>
	0xE642: '襭' // U+896D <cjk>
	0xE643: '襪' // U+896A <cjk>
	0xE644: '襯' // U+896F <cjk>
	0xE645: '襴' // U+8974 <cjk>
	0xE646: '襷' // U+8977 <cjk>
	0xE647: '襾' // U+897E <cjk>
	0xE648: '覃' // U+8983 <cjk>
	0xE649: '覈' // U+8988 <cjk>
	0xE64A: '覊' // U+898A <cjk>
	0xE64B: '覓' // U+8993 <cjk>
	0xE64C: '覘' // U+8998 <cjk>
	0xE64D: '覡' // U+89A1 <cjk>
	0xE64E: '覩' // U+89A9 <cjk>
	0xE64F: '覦' // U+89A6 <cjk>
	0xE650: '覬' // U+89AC <cjk>
	0xE651: '覯' // U+89AF <cjk>
	0xE652: '覲' // U+89B2 <cjk>
	0xE653: '覺' // U+89BA <cjk>
	0xE654: '覽' // U+89BD <cjk>
	0xE655: '覿' // U+89BF <cjk>
	0xE656: '觀' // U+89C0 <cjk>
	0xE657: '觚' // U+89DA <cjk>
	0xE658: '觜' // U+89DC <cjk>
	0xE659: '觝' // U+89DD <cjk>
	0xE65A: '觧' // U+89E7 <cjk>
	0xE65B: '觴' // U+89F4 <cjk>
	0xE65C: '觸' // U+89F8 <cjk>
	0xE65D: '訃' // U+8A03 <cjk>
	0xE65E: '訖' // U+8A16 <cjk>
	0xE65F: '訐' // U+8A10 <cjk>
	0xE660: '訌' // U+8A0C <cjk>
	0xE661: '訛' // U+8A1B <cjk>
	0xE662: '訝' // U+8A1D <cjk>
	0xE663: '訥' // U+8A25 <cjk>
	0xE664: '訶' // U+8A36 <cjk>
	0xE665: '詁' // U+8A41 <cjk>
	0xE666: '詛' // U+8A5B <cjk>
	0xE667: '詒' // U+8A52 <cjk>
	0xE668: '詆' // U+8A46 <cjk>
	0xE669: '詈' // U+8A48 <cjk>
	0xE66A: '詼' // U+8A7C <cjk>
	0xE66B: '詭' // U+8A6D <cjk>
	0xE66C: '詬' // U+8A6C <cjk>
	0xE66D: '詢' // U+8A62 <cjk>
	0xE66E: '誅' // U+8A85 <cjk>
	0xE66F: '誂' // U+8A82 <cjk>
	0xE670: '誄' // U+8A84 <cjk>
	0xE671: '誨' // U+8AA8 <cjk>
	0xE672: '誡' // U+8AA1 <cjk>
	0xE673: '誑' // U+8A91 <cjk>
	0xE674: '誥' // U+8AA5 <cjk>
	0xE675: '誦' // U+8AA6 <cjk>
	0xE676: '誚' // U+8A9A <cjk>
	0xE677: '誣' // U+8AA3 <cjk>
	0xE678: '諄' // U+8AC4 <cjk>
	0xE679: '諍' // U+8ACD <cjk>
	0xE67A: '諂' // U+8AC2 <cjk>
	0xE67B: '諚' // U+8ADA <cjk>
	0xE67C: '諫' // U+8AEB <cjk>
	0xE67D: '諳' // U+8AF3 <cjk>
	0xE67E: '諧' // U+8AE7 <cjk>
	0xE680: '諤' // U+8AE4 <cjk>
	0xE681: '諱' // U+8AF1 <cjk>
	0xE682: '謔' // U+8B14 <cjk>
	0xE683: '諠' // U+8AE0 <cjk>
	0xE684: '諢' // U+8AE2 <cjk>
	0xE685: '諷' // U+8AF7 <cjk>
	0xE686: '諞' // U+8ADE <cjk>
	0xE687: '諛' // U+8ADB <cjk>
	0xE688: '謌' // U+8B0C <cjk>
	0xE689: '謇' // U+8B07 <cjk>
	0xE68A: '謚' // U+8B1A <cjk>
	0xE68B: '諡' // U+8AE1 <cjk>
	0xE68C: '謖' // U+8B16 <cjk>
	0xE68D: '謐' // U+8B10 <cjk>
	0xE68E: '謗' // U+8B17 <cjk>
	0xE68F: '謠' // U+8B20 <cjk>
	0xE690: '謳' // U+8B33 <cjk>
	0xE691: '鞫' // U+97AB <cjk>
	0xE692: '謦' // U+8B26 <cjk>
	0xE693: '謫' // U+8B2B <cjk>
	0xE694: '謾' // U+8B3E <cjk>
	0xE695: '謨' // U+8B28 <cjk>
	0xE696: '譁' // U+8B41 <cjk>
	0xE697: '譌' // U+8B4C <cjk>
	0xE698: '譏' // U+8B4F <cjk>
	0xE699: '譎' // U+8B4E <cjk>
	0xE69A: '證' // U+8B49 <cjk>
	0xE69B: '譖' // U+8B56 <cjk>
	0xE69C: '譛' // U+8B5B <cjk>
	0xE69D: '譚' // U+8B5A <cjk>
	0xE69E: '譫' // U+8B6B <cjk>
	0xE69F: '譟' // U+8B5F <cjk>
	0xE6A0: '譬' // U+8B6C <cjk>
	0xE6A1: '譯' // U+8B6F <cjk>
	0xE6A2: '譴' // U+8B74 <cjk>
	0xE6A3: '譽' // U+8B7D <cjk>
	0xE6A4: '讀' // U+8B80 <cjk>
	0xE6A5: '讌' // U+8B8C <cjk>
	0xE6A6: '讎' // U+8B8E <cjk>
	0xE6A7: '讒' // U+8B92 <cjk>
	0xE6A8: '讓' // U+8B93 <cjk>
	0xE6A9: '讖' // U+8B96 <cjk>
	0xE6AA: '讙' // U+8B99 <cjk>
	0xE6AB: '讚' // U+8B9A <cjk>
	0xE6AC: '谺' // U+8C3A <cjk>
	0xE6AD: '豁' // U+8C41 <cjk>
	0xE6AE: '谿' // U+8C3F <cjk>
	0xE6AF: '豈' // U+8C48 <cjk>
	0xE6B0: '豌' // U+8C4C <cjk>
	0xE6B1: '豎' // U+8C4E <cjk>
	0xE6B2: '豐' // U+8C50 <cjk>
	0xE6B3: '豕' // U+8C55 <cjk>
	0xE6B4: '豢' // U+8C62 <cjk>
	0xE6B5: '豬' // U+8C6C <cjk>
	0xE6B6: '豸' // U+8C78 <cjk>
	0xE6B7: '豺' // U+8C7A <cjk>
	0xE6B8: '貂' // U+8C82 <cjk>
	0xE6B9: '貉' // U+8C89 <cjk>
	0xE6BA: '貅' // U+8C85 <cjk>
	0xE6BB: '貊' // U+8C8A <cjk>
	0xE6BC: '貍' // U+8C8D <cjk>
	0xE6BD: '貎' // U+8C8E <cjk>
	0xE6BE: '貔' // U+8C94 <cjk>
	0xE6BF: '豼' // U+8C7C <cjk>
	0xE6C0: '貘' // U+8C98 <cjk>
	0xE6C1: '戝' // U+621D <cjk>
	0xE6C2: '貭' // U+8CAD <cjk>
	0xE6C3: '貪' // U+8CAA <cjk>
	0xE6C4: '貽' // U+8CBD <cjk>
	0xE6C5: '貲' // U+8CB2 <cjk>
	0xE6C6: '貳' // U+8CB3 <cjk>
	0xE6C7: '貮' // U+8CAE <cjk>
	0xE6C8: '貶' // U+8CB6 <cjk>
	0xE6C9: '賈' // U+8CC8 <cjk>
	0xE6CA: '賁' // U+8CC1 <cjk>
	0xE6CB: '賤' // U+8CE4 <cjk>
	0xE6CC: '賣' // U+8CE3 <cjk>
	0xE6CD: '賚' // U+8CDA <cjk>
	0xE6CE: '賽' // U+8CFD <cjk>
	0xE6CF: '賺' // U+8CFA <cjk>
	0xE6D0: '賻' // U+8CFB <cjk>
	0xE6D1: '贄' // U+8D04 <cjk>
	0xE6D2: '贅' // U+8D05 <cjk>
	0xE6D3: '贊' // U+8D0A <cjk>
	0xE6D4: '贇' // U+8D07 <cjk>
	0xE6D5: '贏' // U+8D0F <cjk>
	0xE6D6: '贍' // U+8D0D <cjk>
	0xE6D7: '贐' // U+8D10 <cjk>
	0xE6D8: '齎' // U+9F4E <cjk>
	0xE6D9: '贓' // U+8D13 <cjk>
	0xE6DA: '賍' // U+8CCD <cjk>
	0xE6DB: '贔' // U+8D14 <cjk>
	0xE6DC: '贖' // U+8D16 <cjk>
	0xE6DD: '赧' // U+8D67 <cjk>
	0xE6DE: '赭' // U+8D6D <cjk>
	0xE6DF: '赱' // U+8D71 <cjk>
	0xE6E0: '赳' // U+8D73 <cjk>
	0xE6E1: '趁' // U+8D81 <cjk>
	0xE6E2: '趙' // U+8D99 <cjk>
	0xE6E3: '跂' // U+8DC2 <cjk>
	0xE6E4: '趾' // U+8DBE <cjk>
	0xE6E5: '趺' // U+8DBA <cjk>
	0xE6E6: '跏' // U+8DCF <cjk>
	0xE6E7: '跚' // U+8DDA <cjk>
	0xE6E8: '跖' // U+8DD6 <cjk>
	0xE6E9: '跌' // U+8DCC <cjk>
	0xE6EA: '跛' // U+8DDB <cjk>
	0xE6EB: '跋' // U+8DCB <cjk>
	0xE6EC: '跪' // U+8DEA <cjk>
	0xE6ED: '跫' // U+8DEB <cjk>
	0xE6EE: '跟' // U+8DDF <cjk>
	0xE6EF: '跣' // U+8DE3 <cjk>
	0xE6F0: '跼' // U+8DFC <cjk>
	0xE6F1: '踈' // U+8E08 <cjk>
	0xE6F2: '踉' // U+8E09 <cjk>
	0xE6F3: '跿' // U+8DFF <cjk>
	0xE6F4: '踝' // U+8E1D <cjk>
	0xE6F5: '踞' // U+8E1E <cjk>
	0xE6F6: '踐' // U+8E10 <cjk>
	0xE6F7: '踟' // U+8E1F <cjk>
	0xE6F8: '蹂' // U+8E42 <cjk>
	0xE6F9: '踵' // U+8E35 <cjk>
	0xE6FA: '踰' // U+8E30 <cjk>
	0xE6FB: '踴' // U+8E34 <cjk>
	0xE6FC: '蹊' // U+8E4A <cjk>
	0xE740: '蹇' // U+8E47 <cjk>
	0xE741: '蹉' // U+8E49 <cjk>
	0xE742: '蹌' // U+8E4C <cjk>
	0xE743: '蹐' // U+8E50 <cjk>
	0xE744: '蹈' // U+8E48 <cjk>
	0xE745: '蹙' // U+8E59 <cjk>
	0xE746: '蹤' // U+8E64 <cjk>
	0xE747: '蹠' // U+8E60 <cjk>
	0xE748: '踪' // U+8E2A <cjk>
	0xE749: '蹣' // U+8E63 <cjk>
	0xE74A: '蹕' // U+8E55 <cjk>
	0xE74B: '蹶' // U+8E76 <cjk>
	0xE74C: '蹲' // U+8E72 <cjk>
	0xE74D: '蹼' // U+8E7C <cjk>
	0xE74E: '躁' // U+8E81 <cjk>
	0xE74F: '躇' // U+8E87 <cjk>
	0xE750: '躅' // U+8E85 <cjk>
	0xE751: '躄' // U+8E84 <cjk>
	0xE752: '躋' // U+8E8B <cjk>
	0xE753: '躊' // U+8E8A <cjk>
	0xE754: '躓' // U+8E93 <cjk>
	0xE755: '躑' // U+8E91 <cjk>
	0xE756: '躔' // U+8E94 <cjk>
	0xE757: '躙' // U+8E99 <cjk>
	0xE758: '躪' // U+8EAA <cjk>
	0xE759: '躡' // U+8EA1 <cjk>
	0xE75A: '躬' // U+8EAC <cjk>
	0xE75B: '躰' // U+8EB0 <cjk>
	0xE75C: '軆' // U+8EC6 <cjk>
	0xE75D: '躱' // U+8EB1 <cjk>
	0xE75E: '躾' // U+8EBE <cjk>
	0xE75F: '軅' // U+8EC5 <cjk>
	0xE760: '軈' // U+8EC8 <cjk>
	0xE761: '軋' // U+8ECB <cjk>
	0xE762: '軛' // U+8EDB <cjk>
	0xE763: '軣' // U+8EE3 <cjk>
	0xE764: '軼' // U+8EFC <cjk>
	0xE765: '軻' // U+8EFB <cjk>
	0xE766: '軫' // U+8EEB <cjk>
	0xE767: '軾' // U+8EFE <cjk>
	0xE768: '輊' // U+8F0A <cjk>
	0xE769: '輅' // U+8F05 <cjk>
	0xE76A: '輕' // U+8F15 <cjk>
	0xE76B: '輒' // U+8F12 <cjk>
	0xE76C: '輙' // U+8F19 <cjk>
	0xE76D: '輓' // U+8F13 <cjk>
	0xE76E: '輜' // U+8F1C <cjk>
	0xE76F: '輟' // U+8F1F <cjk>
	0xE770: '輛' // U+8F1B <cjk>
	0xE771: '輌' // U+8F0C <cjk>
	0xE772: '輦' // U+8F26 <cjk>
	0xE773: '輳' // U+8F33 <cjk>
	0xE774: '輻' // U+8F3B <cjk>
	0xE775: '輹' // U+8F39 <cjk>
	0xE776: '轅' // U+8F45 <cjk>
	0xE777: '轂' // U+8F42 <cjk>
	0xE778: '輾' // U+8F3E <cjk>
	0xE779: '轌' // U+8F4C <cjk>
	0xE77A: '轉' // U+8F49 <cjk>
	0xE77B: '轆' // U+8F46 <cjk>
	0xE77C: '轎' // U+8F4E <cjk>
	0xE77D: '轗' // U+8F57 <cjk>
	0xE77E: '轜' // U+8F5C <cjk>
	0xE780: '轢' // U+8F62 <cjk>
	0xE781: '轣' // U+8F63 <cjk>
	0xE782: '轤' // U+8F64 <cjk>
	0xE783: '辜' // U+8F9C <cjk>
	0xE784: '辟' // U+8F9F <cjk>
	0xE785: '辣' // U+8FA3 <cjk>
	0xE786: '辭' // U+8FAD <cjk>
	0xE787: '辯' // U+8FAF <cjk>
	0xE788: '辷' // U+8FB7 <cjk>
	0xE789: '迚' // U+8FDA <cjk>
	0xE78A: '迥' // U+8FE5 <cjk>
	0xE78B: '迢' // U+8FE2 <cjk>
	0xE78C: '迪' // U+8FEA <cjk>
	0xE78D: '迯' // U+8FEF <cjk>
	0xE78E: '邇' // U+9087 <cjk>
	0xE78F: '迴' // U+8FF4 <cjk>
	0xE790: '逅' // U+9005 <cjk>
	0xE791: '迹' // U+8FF9 <cjk>
	0xE792: '迺' // U+8FFA <cjk>
	0xE793: '逑' // U+9011 <cjk>
	0xE794: '逕' // U+9015 <cjk>
	0xE795: '逡' // U+9021 <cjk>
	0xE796: '逍' // U+900D <cjk>
	0xE797: '逞' // U+901E <cjk>
	0xE798: '逖' // U+9016 <cjk>
	0xE799: '逋' // U+900B <cjk>
	0xE79A: '逧' // U+9027 <cjk>
	0xE79B: '逶' // U+9036 <cjk>
	0xE79C: '逵' // U+9035 <cjk>
	0xE79D: '逹' // U+9039 <cjk>
	0xE79E: '迸' // U+8FF8 <cjk>
	0xE79F: '遏' // U+904F <cjk>
	0xE7A0: '遐' // U+9050 <cjk>
	0xE7A1: '遑' // U+9051 <cjk>
	0xE7A2: '遒' // U+9052 <cjk>
	0xE7A3: '逎' // U+900E <cjk>
	0xE7A4: '遉' // U+9049 <cjk>
	0xE7A5: '逾' // U+903E <cjk>
	0xE7A6: '遖' // U+9056 <cjk>
	0xE7A7: '遘' // U+9058 <cjk>
	0xE7A8: '遞' // U+905E <cjk>
	0xE7A9: '遨' // U+9068 <cjk>
	0xE7AA: '遯' // U+906F <cjk>
	0xE7AB: '遶' // U+9076 <cjk>
	0xE7AC: '隨' // U+96A8 <cjk>
	0xE7AD: '遲' // U+9072 <cjk>
	0xE7AE: '邂' // U+9082 <cjk>
	0xE7AF: '遽' // U+907D <cjk>
	0xE7B0: '邁' // U+9081 <cjk>
	0xE7B1: '邀' // U+9080 <cjk>
	0xE7B2: '邊' // U+908A <cjk>
	0xE7B3: '邉' // U+9089 <cjk>
	0xE7B4: '邏' // U+908F <cjk>
	0xE7B5: '邨' // U+90A8 <cjk>
	0xE7B6: '邯' // U+90AF <cjk>
	0xE7B7: '邱' // U+90B1 <cjk>
	0xE7B8: '邵' // U+90B5 <cjk>
	0xE7B9: '郢' // U+90E2 <cjk>
	0xE7BA: '郤' // U+90E4 <cjk>
	0xE7BB: '扈' // U+6248 <cjk>
	0xE7BC: '郛' // U+90DB <cjk>
	0xE7BD: '鄂' // U+9102 <cjk>
	0xE7BE: '鄒' // U+9112 <cjk>
	0xE7BF: '鄙' // U+9119 <cjk>
	0xE7C0: '鄲' // U+9132 <cjk>
	0xE7C1: '鄰' // U+9130 <cjk>
	0xE7C2: '酊' // U+914A <cjk>
	0xE7C3: '酖' // U+9156 <cjk>
	0xE7C4: '酘' // U+9158 <cjk>
	0xE7C5: '酣' // U+9163 <cjk>
	0xE7C6: '酥' // U+9165 <cjk>
	0xE7C7: '酩' // U+9169 <cjk>
	0xE7C8: '酳' // U+9173 <cjk>
	0xE7C9: '酲' // U+9172 <cjk>
	0xE7CA: '醋' // U+918B <cjk>
	0xE7CB: '醉' // U+9189 <cjk>
	0xE7CC: '醂' // U+9182 <cjk>
	0xE7CD: '醢' // U+91A2 <cjk>
	0xE7CE: '醫' // U+91AB <cjk>
	0xE7CF: '醯' // U+91AF <cjk>
	0xE7D0: '醪' // U+91AA <cjk>
	0xE7D1: '醵' // U+91B5 <cjk>
	0xE7D2: '醴' // U+91B4 <cjk>
	0xE7D3: '醺' // U+91BA <cjk>
	0xE7D4: '釀' // U+91C0 <cjk>
	0xE7D5: '釁' // U+91C1 <cjk>
	0xE7D6: '釉' // U+91C9 <cjk>
	0xE7D7: '釋' // U+91CB <cjk>
	0xE7D8: '釐' // U+91D0 <cjk>
	0xE7D9: '釖' // U+91D6 <cjk>
	0xE7DA: '釟' // U+91DF <cjk>
	0xE7DB: '釡' // U+91E1 <cjk>
	0xE7DC: '釛' // U+91DB <cjk>
	0xE7DD: '釼' // U+91FC <cjk>
	0xE7DE: '釵' // U+91F5 <cjk>
	0xE7DF: '釶' // U+91F6 <cjk>
	0xE7E0: '鈞' // U+921E <cjk>
	0xE7E1: '釿' // U+91FF <cjk>
	0xE7E2: '鈔' // U+9214 <cjk>
	0xE7E3: '鈬' // U+922C <cjk>
	0xE7E4: '鈕' // U+9215 <cjk>
	0xE7E5: '鈑' // U+9211 <cjk>
	0xE7E6: '鉞' // U+925E <cjk>
	0xE7E7: '鉗' // U+9257 <cjk>
	0xE7E8: '鉅' // U+9245 <cjk>
	0xE7E9: '鉉' // U+9249 <cjk>
	0xE7EA: '鉤' // U+9264 <cjk>
	0xE7EB: '鉈' // U+9248 <cjk>
	0xE7EC: '銕' // U+9295 <cjk>
	0xE7ED: '鈿' // U+923F <cjk>
	0xE7EE: '鉋' // U+924B <cjk>
	0xE7EF: '鉐' // U+9250 <cjk>
	0xE7F0: '銜' // U+929C <cjk>
	0xE7F1: '銖' // U+9296 <cjk>
	0xE7F2: '銓' // U+9293 <cjk>
	0xE7F3: '銛' // U+929B <cjk>
	0xE7F4: '鉚' // U+925A <cjk>
	0xE7F5: '鋏' // U+92CF <cjk>
	0xE7F6: '銹' // U+92B9 <cjk>
	0xE7F7: '銷' // U+92B7 <cjk>
	0xE7F8: '鋩' // U+92E9 <cjk>
	0xE7F9: '錏' // U+930F <cjk>
	0xE7FA: '鋺' // U+92FA <cjk>
	0xE7FB: '鍄' // U+9344 <cjk>
	0xE7FC: '錮' // U+932E <cjk>
	0xE840: '錙' // U+9319 <cjk>
	0xE841: '錢' // U+9322 <cjk>
	0xE842: '錚' // U+931A <cjk>
	0xE843: '錣' // U+9323 <cjk>
	0xE844: '錺' // U+933A <cjk>
	0xE845: '錵' // U+9335 <cjk>
	0xE846: '錻' // U+933B <cjk>
	0xE847: '鍜' // U+935C <cjk>
	0xE848: '鍠' // U+9360 <cjk>
	0xE849: '鍼' // U+937C <cjk>
	0xE84A: '鍮' // U+936E <cjk>
	0xE84B: '鍖' // U+9356 <cjk>
	0xE84C: '鎰' // U+93B0 <cjk>
	0xE84D: '鎬' // U+93AC <cjk>
	0xE84E: '鎭' // U+93AD <cjk>
	0xE84F: '鎔' // U+9394 <cjk>
	0xE850: '鎹' // U+93B9 <cjk>
	0xE851: '鏖' // U+93D6 <cjk>
	0xE852: '鏗' // U+93D7 <cjk>
	0xE853: '鏨' // U+93E8 <cjk>
	0xE854: '鏥' // U+93E5 <cjk>
	0xE855: '鏘' // U+93D8 <cjk>
	0xE856: '鏃' // U+93C3 <cjk>
	0xE857: '鏝' // U+93DD <cjk>
	0xE858: '鏐' // U+93D0 <cjk>
	0xE859: '鏈' // U+93C8 <cjk>
	0xE85A: '鏤' // U+93E4 <cjk>
	0xE85B: '鐚' // U+941A <cjk>
	0xE85C: '鐔' // U+9414 <cjk>
	0xE85D: '鐓' // U+9413 <cjk>
	0xE85E: '鐃' // U+9403 <cjk>
	0xE85F: '鐇' // U+9407 <cjk>
	0xE860: '鐐' // U+9410 <cjk>
	0xE861: '鐶' // U+9436 <cjk>
	0xE862: '鐫' // U+942B <cjk>
	0xE863: '鐵' // U+9435 <cjk>
	0xE864: '鐡' // U+9421 <cjk>
	0xE865: '鐺' // U+943A <cjk>
	0xE866: '鑁' // U+9441 <cjk>
	0xE867: '鑒' // U+9452 <cjk>
	0xE868: '鑄' // U+9444 <cjk>
	0xE869: '鑛' // U+945B <cjk>
	0xE86A: '鑠' // U+9460 <cjk>
	0xE86B: '鑢' // U+9462 <cjk>
	0xE86C: '鑞' // U+945E <cjk>
	0xE86D: '鑪' // U+946A <cjk>
	0xE86E: '鈩' // U+9229 <cjk>
	0xE86F: '鑰' // U+9470 <cjk>
	0xE870: '鑵' // U+9475 <cjk>
	0xE871: '鑷' // U+9477 <cjk>
	0xE872: '鑽' // U+947D <cjk>
	0xE873: '鑚' // U+945A <cjk>
	0xE874: '鑼' // U+947C <cjk>
	0xE875: '鑾' // U+947E <cjk>
	0xE876: '钁' // U+9481 <cjk>
	0xE877: '鑿' // U+947F <cjk>
	0xE878: '閂' // U+9582 <cjk>
	0xE879: '閇' // U+9587 <cjk>
	0xE87A: '閊' // U+958A <cjk>
	0xE87B: '閔' // U+9594 <cjk>
	0xE87C: '閖' // U+9596 <cjk>
	0xE87D: '閘' // U+9598 <cjk>
	0xE87E: '閙' // U+9599 <cjk>
	0xE880: '閠' // U+95A0 <cjk>
	0xE881: '閨' // U+95A8 <cjk>
	0xE882: '閧' // U+95A7 <cjk>
	0xE883: '閭' // U+95AD <cjk>
	0xE884: '閼' // U+95BC <cjk>
	0xE885: '閻' // U+95BB <cjk>
	0xE886: '閹' // U+95B9 <cjk>
	0xE887: '閾' // U+95BE <cjk>
	0xE888: '闊' // U+95CA <cjk>
	0xE889: '濶' // U+6FF6 <cjk>
	0xE88A: '闃' // U+95C3 <cjk>
	0xE88B: '闍' // U+95CD <cjk>
	0xE88C: '闌' // U+95CC <cjk>
	0xE88D: '闕' // U+95D5 <cjk>
	0xE88E: '闔' // U+95D4 <cjk>
	0xE88F: '闖' // U+95D6 <cjk>
	0xE890: '關' // U+95DC <cjk>
	0xE891: '闡' // U+95E1 <cjk>
	0xE892: '闥' // U+95E5 <cjk>
	0xE893: '闢' // U+95E2 <cjk>
	0xE894: '阡' // U+9621 <cjk>
	0xE895: '阨' // U+9628 <cjk>
	0xE896: '阮' // U+962E <cjk>
	0xE897: '阯' // U+962F <cjk>
	0xE898: '陂' // U+9642 <cjk>
	0xE899: '陌' // U+964C <cjk>
	0xE89A: '陏' // U+964F <cjk>
	0xE89B: '陋' // U+964B <cjk>
	0xE89C: '陷' // U+9677 <cjk>
	0xE89D: '陜' // U+965C <cjk>
	0xE89E: '陞' // U+965E <cjk>
	0xE89F: '陝' // U+965D <cjk>
	0xE8A0: '陟' // U+965F <cjk>
	0xE8A1: '陦' // U+9666 <cjk>
	0xE8A2: '陲' // U+9672 <cjk>
	0xE8A3: '陬' // U+966C <cjk>
	0xE8A4: '隍' // U+968D <cjk>
	0xE8A5: '隘' // U+9698 <cjk>
	0xE8A6: '隕' // U+9695 <cjk>
	0xE8A7: '隗' // U+9697 <cjk>
	0xE8A8: '險' // U+96AA <cjk>
	0xE8A9: '隧' // U+96A7 <cjk>
	0xE8AA: '隱' // U+96B1 <cjk>
	0xE8AB: '隲' // U+96B2 <cjk>
	0xE8AC: '隰' // U+96B0 <cjk>
	0xE8AD: '隴' // U+96B4 <cjk>
	0xE8AE: '隶' // U+96B6 <cjk>
	0xE8AF: '隸' // U+96B8 <cjk>
	0xE8B0: '隹' // U+96B9 <cjk>
	0xE8B1: '雎' // U+96CE <cjk>
	0xE8B2: '雋' // U+96CB <cjk>
	0xE8B3: '雉' // U+96C9 <cjk>
	0xE8B4: '雍' // U+96CD <cjk>
	0xE8B5: '襍' // U+894D <cjk>
	0xE8B6: '雜' // U+96DC <cjk>
	0xE8B7: '霍' // U+970D <cjk>
	0xE8B8: '雕' // U+96D5 <cjk>
	0xE8B9: '雹' // U+96F9 <cjk>
	0xE8BA: '霄' // U+9704 <cjk>
	0xE8BB: '霆' // U+9706 <cjk>
	0xE8BC: '霈' // U+9708 <cjk>
	0xE8BD: '霓' // U+9713 <cjk>
	0xE8BE: '霎' // U+970E <cjk>
	0xE8BF: '霑' // U+9711 <cjk>
	0xE8C0: '霏' // U+970F <cjk>
	0xE8C1: '霖' // U+9716 <cjk>
	0xE8C2: '霙' // U+9719 <cjk>
	0xE8C3: '霤' // U+9724 <cjk>
	0xE8C4: '霪' // U+972A <cjk>
	0xE8C5: '霰' // U+9730 <cjk>
	0xE8C6: '霹' // U+9739 <cjk>
	0xE8C7: '霽' // U+973D <cjk>
	0xE8C8: '霾' // U+973E <cjk>
	0xE8C9: '靄' // U+9744 <cjk>
	0xE8CA: '靆' // U+9746 <cjk>
	0xE8CB: '靈' // U+9748 <cjk>
	0xE8CC: '靂' // U+9742 <cjk>
	0xE8CD: '靉' // U+9749 <cjk>
	0xE8CE: '靜' // U+975C <cjk>
	0xE8CF: '靠' // U+9760 <cjk>
	0xE8D0: '靤' // U+9764 <cjk>
	0xE8D1: '靦' // U+9766 <cjk>
	0xE8D2: '靨' // U+9768 <cjk>
	0xE8D3: '勒' // U+52D2 <cjk>
	0xE8D4: '靫' // U+976B <cjk>
	0xE8D5: '靱' // U+9771 <cjk>
	0xE8D6: '靹' // U+9779 <cjk>
	0xE8D7: '鞅' // U+9785 <cjk>
	0xE8D8: '靼' // U+977C <cjk>
	0xE8D9: '鞁' // U+9781 <cjk>
	0xE8DA: '靺' // U+977A <cjk>
	0xE8DB: '鞆' // U+9786 <cjk>
	0xE8DC: '鞋' // U+978B <cjk>
	0xE8DD: '鞏' // U+978F <cjk>
	0xE8DE: '鞐' // U+9790 <cjk>
	0xE8DF: '鞜' // U+979C <cjk>
	0xE8E0: '鞨' // U+97A8 <cjk>
	0xE8E1: '鞦' // U+97A6 <cjk>
	0xE8E2: '鞣' // U+97A3 <cjk>
	0xE8E3: '鞳' // U+97B3 <cjk>
	0xE8E4: '鞴' // U+97B4 <cjk>
	0xE8E5: '韃' // U+97C3 <cjk>
	0xE8E6: '韆' // U+97C6 <cjk>
	0xE8E7: '韈' // U+97C8 <cjk>
	0xE8E8: '韋' // U+97CB <cjk>
	0xE8E9: '韜' // U+97DC <cjk>
	0xE8EA: '韭' // U+97ED <cjk>
	0xE8EB: '齏' // U+9F4F <cjk>
	0xE8EC: '韲' // U+97F2 <cjk>
	0xE8ED: '竟' // U+7ADF <cjk>
	0xE8EE: '韶' // U+97F6 <cjk>
	0xE8EF: '韵' // U+97F5 <cjk>
	0xE8F0: '頏' // U+980F <cjk>
	0xE8F1: '頌' // U+980C <cjk>
	0xE8F2: '頸' // U+9838 <cjk>
	0xE8F3: '頤' // U+9824 <cjk>
	0xE8F4: '頡' // U+9821 <cjk>
	0xE8F5: '頷' // U+9837 <cjk>
	0xE8F6: '頽' // U+983D <cjk>
	0xE8F7: '顆' // U+9846 <cjk>
	0xE8F8: '顏' // U+984F <cjk>
	0xE8F9: '顋' // U+984B <cjk>
	0xE8FA: '顫' // U+986B <cjk>
	0xE8FB: '顯' // U+986F <cjk>
	0xE8FC: '顰' // U+9870 <cjk>
	0xE940: '顱' // U+9871 <cjk>
	0xE941: '顴' // U+9874 <cjk>
	0xE942: '顳' // U+9873 <cjk>
	0xE943: '颪' // U+98AA <cjk>
	0xE944: '颯' // U+98AF <cjk>
	0xE945: '颱' // U+98B1 <cjk>
	0xE946: '颶' // U+98B6 <cjk>
	0xE947: '飄' // U+98C4 <cjk>
	0xE948: '飃' // U+98C3 <cjk>
	0xE949: '飆' // U+98C6 <cjk>
	0xE94A: '飩' // U+98E9 <cjk>
	0xE94B: '飫' // U+98EB <cjk>
	0xE94C: '餃' // U+9903 <cjk>
	0xE94D: '餉' // U+9909 <cjk>
	0xE94E: '餒' // U+9912 <cjk>
	0xE94F: '餔' // U+9914 <cjk>
	0xE950: '餘' // U+9918 <cjk>
	0xE951: '餡' // U+9921 <cjk>
	0xE952: '餝' // U+991D <cjk>
	0xE953: '餞' // U+991E <cjk>
	0xE954: '餤' // U+9924 <cjk>
	0xE955: '餠' // U+9920 <cjk>
	0xE956: '餬' // U+992C <cjk>
	0xE957: '餮' // U+992E <cjk>
	0xE958: '餽' // U+993D <cjk>
	0xE959: '餾' // U+993E <cjk>
	0xE95A: '饂' // U+9942 <cjk>
	0xE95B: '饉' // U+9949 <cjk>
	0xE95C: '饅' // U+9945 <cjk>
	0xE95D: '饐' // U+9950 <cjk>
	0xE95E: '饋' // U+994B <cjk>
	0xE95F: '饑' // U+9951 <cjk>
	0xE960: '饒' // U+9952 <cjk>
	0xE961: '饌' // U+994C <cjk>
	0xE962: '饕' // U+9955 <cjk>
	0xE963: '馗' // U+9997 <cjk>
	0xE964: '馘' // U+9998 <cjk>
	0xE965: '馥' // U+99A5 <cjk>
	0xE966: '馭' // U+99AD <cjk>
	0xE967: '馮' // U+99AE <cjk>
	0xE968: '馼' // U+99BC <cjk>
	0xE969: '駟' // U+99DF <cjk>
	0xE96A: '駛' // U+99DB <cjk>
	0xE96B: '駝' // U+99DD <cjk>
	0xE96C: '駘' // U+99D8 <cjk>
	0xE96D: '駑' // U+99D1 <cjk>
	0xE96E: '駭' // U+99ED <cjk>
	0xE96F: '駮' // U+99EE <cjk>
	0xE970: '駱' // U+99F1 <cjk>
	0xE971: '駲' // U+99F2 <cjk>
	0xE972: '駻' // U+99FB <cjk>
	0xE973: '駸' // U+99F8 <cjk>
	0xE974: '騁' // U+9A01 <cjk>
	0xE975: '騏' // U+9A0F <cjk>
	0xE976: '騅' // U+9A05 <cjk>
	0xE977: '駢' // U+99E2 <cjk>
	0xE978: '騙' // U+9A19 <cjk>
	0xE979: '騫' // U+9A2B <cjk>
	0xE97A: '騷' // U+9A37 <cjk>
	0xE97B: '驅' // U+9A45 <cjk>
	0xE97C: '驂' // U+9A42 <cjk>
	0xE97D: '驀' // U+9A40 <cjk>
	0xE97E: '驃' // U+9A43 <cjk>
	0xE980: '騾' // U+9A3E <cjk>
	0xE981: '驕' // U+9A55 <cjk>
	0xE982: '驍' // U+9A4D <cjk>
	0xE983: '驛' // U+9A5B <cjk>
	0xE984: '驗' // U+9A57 <cjk>
	0xE985: '驟' // U+9A5F <cjk>
	0xE986: '驢' // U+9A62 <cjk>
	0xE987: '驥' // U+9A65 <cjk>
	0xE988: '驤' // U+9A64 <cjk>
	0xE989: '驩' // U+9A69 <cjk>
	0xE98A: '驫' // U+9A6B <cjk>
	0xE98B: '驪' // U+9A6A <cjk>
	0xE98C: '骭' // U+9AAD <cjk>
	0xE98D: '骰' // U+9AB0 <cjk>
	0xE98E: '骼' // U+9ABC <cjk>
	0xE98F: '髀' // U+9AC0 <cjk>
	0xE990: '髏' // U+9ACF <cjk>
	0xE991: '髑' // U+9AD1 <cjk>
	0xE992: '髓' // U+9AD3 <cjk>
	0xE993: '體' // U+9AD4 <cjk>
	0xE994: '髞' // U+9ADE <cjk>
	0xE995: '髟' // U+9ADF <cjk>
	0xE996: '髢' // U+9AE2 <cjk>
	0xE997: '髣' // U+9AE3 <cjk>
	0xE998: '髦' // U+9AE6 <cjk>
	0xE999: '髯' // U+9AEF <cjk>
	0xE99A: '髫' // U+9AEB <cjk>
	0xE99B: '髮' // U+9AEE <cjk>
	0xE99C: '髴' // U+9AF4 <cjk>
	0xE99D: '髱' // U+9AF1 <cjk>
	0xE99E: '髷' // U+9AF7 <cjk>
	0xE99F: '髻' // U+9AFB <cjk>
	0xE9A0: '鬆' // U+9B06 <cjk>
	0xE9A1: '鬘' // U+9B18 <cjk>
	0xE9A2: '鬚' // U+9B1A <cjk>
	0xE9A3: '鬟' // U+9B1F <cjk>
	0xE9A4: '鬢' // U+9B22 <cjk>
	0xE9A5: '鬣' // U+9B23 <cjk>
	0xE9A6: '鬥' // U+9B25 <cjk>
	0xE9A7: '鬧' // U+9B27 <cjk>
	0xE9A8: '鬨' // U+9B28 <cjk>
	0xE9A9: '鬩' // U+9B29 <cjk>
	0xE9AA: '鬪' // U+9B2A <cjk>
	0xE9AB: '鬮' // U+9B2E <cjk>
	0xE9AC: '鬯' // U+9B2F <cjk>
	0xE9AD: '鬲' // U+9B32 <cjk>
	0xE9AE: '魄' // U+9B44 <cjk>
	0xE9AF: '魃' // U+9B43 <cjk>
	0xE9B0: '魏' // U+9B4F <cjk>
	0xE9B1: '魍' // U+9B4D <cjk>
	0xE9B2: '魎' // U+9B4E <cjk>
	0xE9B3: '魑' // U+9B51 <cjk>
	0xE9B4: '魘' // U+9B58 <cjk>
	0xE9B5: '魴' // U+9B74 <cjk>
	0xE9B6: '鮓' // U+9B93 <cjk>
	0xE9B7: '鮃' // U+9B83 <cjk>
	0xE9B8: '鮑' // U+9B91 <cjk>
	0xE9B9: '鮖' // U+9B96 <cjk>
	0xE9BA: '鮗' // U+9B97 <cjk>
	0xE9BB: '鮟' // U+9B9F <cjk>
	0xE9BC: '鮠' // U+9BA0 <cjk>
	0xE9BD: '鮨' // U+9BA8 <cjk>
	0xE9BE: '鮴' // U+9BB4 <cjk>
	0xE9BF: '鯀' // U+9BC0 <cjk>
	0xE9C0: '鯊' // U+9BCA <cjk>
	0xE9C1: '鮹' // U+9BB9 <cjk>
	0xE9C2: '鯆' // U+9BC6 <cjk>
	0xE9C3: '鯏' // U+9BCF <cjk>
	0xE9C4: '鯑' // U+9BD1 <cjk>
	0xE9C5: '鯒' // U+9BD2 <cjk>
	0xE9C6: '鯣' // U+9BE3 <cjk>
	0xE9C7: '鯢' // U+9BE2 <cjk>
	0xE9C8: '鯤' // U+9BE4 <cjk>
	0xE9C9: '鯔' // U+9BD4 <cjk>
	0xE9CA: '鯡' // U+9BE1 <cjk>
	0xE9CB: '鰺' // U+9C3A <cjk>
	0xE9CC: '鯲' // U+9BF2 <cjk>
	0xE9CD: '鯱' // U+9BF1 <cjk>
	0xE9CE: '鯰' // U+9BF0 <cjk>
	0xE9CF: '鰕' // U+9C15 <cjk>
	0xE9D0: '鰔' // U+9C14 <cjk>
	0xE9D1: '鰉' // U+9C09 <cjk>
	0xE9D2: '鰓' // U+9C13 <cjk>
	0xE9D3: '鰌' // U+9C0C <cjk>
	0xE9D4: '鰆' // U+9C06 <cjk>
	0xE9D5: '鰈' // U+9C08 <cjk>
	0xE9D6: '鰒' // U+9C12 <cjk>
	0xE9D7: '鰊' // U+9C0A <cjk>
	0xE9D8: '鰄' // U+9C04 <cjk>
	0xE9D9: '鰮' // U+9C2E <cjk>
	0xE9DA: '鰛' // U+9C1B <cjk>
	0xE9DB: '鰥' // U+9C25 <cjk>
	0xE9DC: '鰤' // U+9C24 <cjk>
	0xE9DD: '鰡' // U+9C21 <cjk>
	0xE9DE: '鰰' // U+9C30 <cjk>
	0xE9DF: '鱇' // U+9C47 <cjk>
	0xE9E0: '鰲' // U+9C32 <cjk>
	0xE9E1: '鱆' // U+9C46 <cjk>
	0xE9E2: '鰾' // U+9C3E <cjk>
	0xE9E3: '鱚' // U+9C5A <cjk>
	0xE9E4: '鱠' // U+9C60 <cjk>
	0xE9E5: '鱧' // U+9C67 <cjk>
	0xE9E6: '鱶' // U+9C76 <cjk>
	0xE9E7: '鱸' // U+9C78 <cjk>
	0xE9E8: '鳧' // U+9CE7 <cjk>
	0xE9E9: '鳬' // U+9CEC <cjk>
	0xE9EA: '鳰' // U+9CF0 <cjk>
	0xE9EB: '鴉' // U+9D09 <cjk>
	0xE9EC: '鴈' // U+9D08 <cjk>
	0xE9ED: '鳫' // U+9CEB <cjk>
	0xE9EE: '鴃' // U+9D03 <cjk>
	0xE9EF: '鴆' // U+9D06 <cjk>
	0xE9F0: '鴪' // U+9D2A <cjk>
	0xE9F1: '鴦' // U+9D26 <cjk>
	0xE9F2: '鶯' // U+9DAF <cjk>
	0xE9F3: '鴣' // U+9D23 <cjk>
	0xE9F4: '鴟' // U+9D1F <cjk>
	0xE9F5: '鵄' // U+9D44 <cjk>
	0xE9F6: '鴕' // U+9D15 <cjk>
	0xE9F7: '鴒' // U+9D12 <cjk>
	0xE9F8: '鵁' // U+9D41 <cjk>
	0xE9F9: '鴿' // U+9D3F <cjk>
	0xE9FA: '鴾' // U+9D3E <cjk>
	0xE9FB: '鵆' // U+9D46 <cjk>
	0xE9FC: '鵈' // U+9D48 <cjk>
	0xEA40: '鵝' // U+9D5D <cjk>
	0xEA41: '鵞' // U+9D5E <cjk>
	0xEA42: '鵤' // U+9D64 <cjk>
	0xEA43: '鵑' // U+9D51 <cjk>
	0xEA44: '鵐' // U+9D50 <cjk>
	0xEA45: '鵙' // U+9D59 <cjk>
	0xEA46: '鵲' // U+9D72 <cjk>
	0xEA47: '鶉' // U+9D89 <cjk>
	0xEA48: '鶇' // U+9D87 <cjk>
	0xEA49: '鶫' // U+9DAB <cjk>
	0xEA4A: '鵯' // U+9D6F <cjk>
	0xEA4B: '鵺' // U+9D7A <cjk>
	0xEA4C: '鶚' // U+9D9A <cjk>
	0xEA4D: '鶤' // U+9DA4 <cjk>
	0xEA4E: '鶩' // U+9DA9 <cjk>
	0xEA4F: '鶲' // U+9DB2 <cjk>
	0xEA50: '鷄' // U+9DC4 <cjk>
	0xEA51: '鷁' // U+9DC1 <cjk>
	0xEA52: '鶻' // U+9DBB <cjk>
	0xEA53: '鶸' // U+9DB8 <cjk>
	0xEA54: '鶺' // U+9DBA <cjk>
	0xEA55: '鷆' // U+9DC6 <cjk>
	0xEA56: '鷏' // U+9DCF <cjk>
	0xEA57: '鷂' // U+9DC2 <cjk>
	0xEA58: '鷙' // U+9DD9 <cjk>
	0xEA59: '鷓' // U+9DD3 <cjk>
	0xEA5A: '鷸' // U+9DF8 <cjk>
	0xEA5B: '鷦' // U+9DE6 <cjk>
	0xEA5C: '鷭' // U+9DED <cjk>
	0xEA5D: '鷯' // U+9DEF <cjk>
	0xEA5E: '鷽' // U+9DFD <cjk>
	0xEA5F: '鸚' // U+9E1A <cjk>
	0xEA60: '鸛' // U+9E1B <cjk>
	0xEA61: '鸞' // U+9E1E <cjk>
	0xEA62: '鹵' // U+9E75 <cjk>
	0xEA63: '鹹' // U+9E79 <cjk>
	0xEA64: '鹽' // U+9E7D <cjk>
	0xEA65: '麁' // U+9E81 <cjk>
	0xEA66: '麈' // U+9E88 <cjk>
	0xEA67: '麋' // U+9E8B <cjk>
	0xEA68: '麌' // U+9E8C <cjk>
	0xEA69: '麒' // U+9E92 <cjk>
	0xEA6A: '麕' // U+9E95 <cjk>
	0xEA6B: '麑' // U+9E91 <cjk>
	0xEA6C: '麝' // U+9E9D <cjk>
	0xEA6D: '麥' // U+9EA5 <cjk>
	0xEA6E: '麩' // U+9EA9 <cjk>
	0xEA6F: '麸' // U+9EB8 <cjk>
	0xEA70: '麪' // U+9EAA <cjk>
	0xEA71: '麭' // U+9EAD <cjk>
	0xEA72: '靡' // U+9761 <cjk>
	0xEA73: '黌' // U+9ECC <cjk>
	0xEA74: '黎' // U+9ECE <cjk>
	0xEA75: '黏' // U+9ECF <cjk>
	0xEA76: '黐' // U+9ED0 <cjk>
	0xEA77: '黔' // U+9ED4 <cjk>
	0xEA78: '黜' // U+9EDC <cjk>
	0xEA79: '點' // U+9EDE <cjk>
	0xEA7A: '黝' // U+9EDD <cjk>
	0xEA7B: '黠' // U+9EE0 <cjk>
	0xEA7C: '黥' // U+9EE5 <cjk>
	0xEA7D: '黨' // U+9EE8 <cjk>
	0xEA7E: '黯' // U+9EEF <cjk>
	0xEA80: '黴' // U+9EF4 <cjk>
	0xEA81: '黶' // U+9EF6 <cjk>
	0xEA82: '黷' // U+9EF7 <cjk>
	0xEA83: '黹' // U+9EF9 <cjk>
	0xEA84: '黻' // U+9EFB <cjk>
	0xEA85: '黼' // U+9EFC <cjk>
	0xEA86: '黽' // U+9EFD <cjk>
	0xEA87: '鼇' // U+9F07 <cjk>
	0xEA88: '鼈' // U+9F08 <cjk>
	0xEA89: '皷' // U+76B7 <cjk>
	0xEA8A: '鼕' // U+9F15 <cjk>
	0xEA8B: '鼡' // U+9F21 <cjk>
	0xEA8C: '鼬' // U+9F2C <cjk>
	0xEA8D: '鼾' // U+9F3E <cjk>
	0xEA8E: '齊' // U+9F4A <cjk>
	0xEA8F: '齒' // U+9F52 <cjk>
	0xEA90: '齔' // U+9F54 <cjk>
	0xEA91: '齣' // U+9F63 <cjk>
	0xEA92: '齟' // U+9F5F <cjk>
	0xEA93: '齠' // U+9F60 <cjk>
	0xEA94: '齡' // U+9F61 <cjk>
	0xEA95: '齦' // U+9F66 <cjk>
	0xEA96: '齧' // U+9F67 <cjk>
	0xEA97: '齬' // U+9F6C <cjk>
	0xEA98: '齪' // U+9F6A <cjk>
	0xEA99: '齷' // U+9F77 <cjk>
	0xEA9A: '齲' // U+9F72 <cjk>
	0xEA9B: '齶' // U+9F76 <cjk>
	0xEA9C: '龕' // U+9F95 <cjk>
	0xEA9D: '龜' // U+9F9C <cjk>
	0xEA9E: '龠' // U+9FA0 <cjk>
	0xEA9F: '堯' // U+582F <cjk>
	0xEAA0: '槇' // U+69C7 <cjk>
	0xEAA1: '遙' // U+9059 <cjk>
	0xEAA2: '瑤' // U+7464 <cjk>
	0xEAA3: '凜' // U+51DC <cjk>
	0xEAA4: '熙' // U+7199 <cjk>
	0xEAA5: '噓' // U+5653 <cjk>
	0xEAA6: '巢' // U+5DE2 <cjk>
	0xEAA7: '帔' // U+5E14 <cjk>
	0xEAA8: '帘' // U+5E18 <cjk>
	0xEAA9: '幘' // U+5E58 <cjk>
	0xEAAA: '幞' // U+5E5E <cjk>
	0xEAAB: '庾' // U+5EBE <cjk>
	0xEAAC: '廊' // U+F928 CJK COMPATIBILITY IDEOGRAPH-F928
	0xEAAD: '廋' // U+5ECB <cjk>
	0xEAAE: '廹' // U+5EF9 <cjk>
	0xEAAF: '开' // U+5F00 <cjk>
	0xEAB0: '异' // U+5F02 <cjk>
	0xEAB1: '弇' // U+5F07 <cjk>
	0xEAB2: '弝' // U+5F1D <cjk>
	0xEAB3: '弣' // U+5F23 <cjk>
	0xEAB4: '弴' // U+5F34 <cjk>
	0xEAB5: '弶' // U+5F36 <cjk>
	0xEAB6: '弽' // U+5F3D <cjk>
	0xEAB7: '彀' // U+5F40 <cjk>
	0xEAB8: '彅' // U+5F45 <cjk>
	0xEAB9: '彔' // U+5F54 <cjk>
	0xEABA: '彘' // U+5F58 <cjk>
	0xEABB: '彤' // U+5F64 <cjk>
	0xEABC: '彧' // U+5F67 <cjk>
	0xEABD: '彽' // U+5F7D <cjk>
	0xEABE: '徉' // U+5F89 <cjk>
	0xEABF: '徜' // U+5F9C <cjk>
	0xEAC0: '徧' // U+5FA7 <cjk>
	0xEAC1: '徯' // U+5FAF <cjk>
	0xEAC2: '徵' // U+5FB5 <cjk>
	0xEAC3: '德' // U+5FB7 <cjk>
	0xEAC4: '忉' // U+5FC9 <cjk>
	0xEAC5: '忞' // U+5FDE <cjk>
	0xEAC6: '忡' // U+5FE1 <cjk>
	0xEAC7: '忩' // U+5FE9 <cjk>
	0xEAC8: '怍' // U+600D <cjk>
	0xEAC9: '怔' // U+6014 <cjk>
	0xEACA: '怘' // U+6018 <cjk>
	0xEACB: '怳' // U+6033 <cjk>
	0xEACC: '怵' // U+6035 <cjk>
	0xEACD: '恇' // U+6047 <cjk>
	0xEACE: '悔' // U+FA3D CJK COMPATIBILITY IDEOGRAPH-FA3D
	0xEACF: '悝' // U+609D <cjk>
	0xEAD0: '悞' // U+609E <cjk>
	0xEAD1: '惋' // U+60CB <cjk>
	0xEAD2: '惔' // U+60D4 <cjk>
	0xEAD3: '惕' // U+60D5 <cjk>
	0xEAD4: '惝' // U+60DD <cjk>
	0xEAD5: '惸' // U+60F8 <cjk>
	0xEAD6: '愜' // U+611C <cjk>
	0xEAD7: '愫' // U+612B <cjk>
	0xEAD8: '愰' // U+6130 <cjk>
	0xEAD9: '愷' // U+6137 <cjk>
	0xEADA: '慨' // U+FA3E CJK COMPATIBILITY IDEOGRAPH-FA3E
	0xEADB: '憍' // U+618D <cjk>
	0xEADC: '憎' // U+FA3F CJK COMPATIBILITY IDEOGRAPH-FA3F
	0xEADD: '憼' // U+61BC <cjk>
	0xEADE: '憹' // U+61B9 <cjk>
	0xEADF: '懲' // U+FA40 CJK COMPATIBILITY IDEOGRAPH-FA40
	0xEAE0: '戢' // U+6222 <cjk>
	0xEAE1: '戾' // U+623E <cjk>
	0xEAE2: '扃' // U+6243 <cjk>
	0xEAE3: '扖' // U+6256 <cjk>
	0xEAE4: '扚' // U+625A <cjk>
	0xEAE5: '扯' // U+626F <cjk>
	0xEAE6: '抅' // U+6285 <cjk>
	0xEAE7: '拄' // U+62C4 <cjk>
	0xEAE8: '拖' // U+62D6 <cjk>
	0xEAE9: '拼' // U+62FC <cjk>
	0xEAEA: '挊' // U+630A <cjk>
	0xEAEB: '挘' // U+6318 <cjk>
	0xEAEC: '挹' // U+6339 <cjk>
	0xEAED: '捃' // U+6343 <cjk>
	0xEAEE: '捥' // U+6365 <cjk>
	0xEAEF: '捼' // U+637C <cjk>
	0xEAF0: '揥' // U+63E5 <cjk>
	0xEAF1: '揭' // U+63ED <cjk>
	0xEAF2: '揵' // U+63F5 <cjk>
	0xEAF3: '搐' // U+6410 <cjk>
	0xEAF4: '搔' // U+6414 <cjk>
	0xEAF5: '搢' // U+6422 <cjk>
	0xEAF6: '摹' // U+6479 <cjk>
	0xEAF7: '摑' // U+6451 <cjk>
	0xEAF8: '摠' // U+6460 <cjk>
	0xEAF9: '摭' // U+646D <cjk>
	0xEAFA: '擎' // U+64CE <cjk>
	0xEAFB: '撾' // U+64BE <cjk>
	0xEAFC: '撿' // U+64BF <cjk>
	0xEB40: '擄' // U+64C4 <cjk>
	0xEB41: '擊' // U+64CA <cjk>
	0xEB42: '擐' // U+64D0 <cjk>
	0xEB43: '擷' // U+64F7 <cjk>
	0xEB44: '擻' // U+64FB <cjk>
	0xEB45: '攢' // U+6522 <cjk>
	0xEB46: '攩' // U+6529 <cjk>
	0xEB47: '敏' // U+FA41 CJK COMPATIBILITY IDEOGRAPH-FA41
	0xEB48: '敧' // U+6567 <cjk>
	0xEB49: '斝' // U+659D <cjk>
	0xEB4A: '既' // U+FA42 CJK COMPATIBILITY IDEOGRAPH-FA42
	0xEB4B: '昀' // U+6600 <cjk>
	0xEB4C: '昉' // U+6609 <cjk>
	0xEB4D: '昕' // U+6615 <cjk>
	0xEB4E: '昞' // U+661E <cjk>
	0xEB4F: '昺' // U+663A <cjk>
	0xEB50: '昢' // U+6622 <cjk>
	0xEB51: '昤' // U+6624 <cjk>
	0xEB52: '昫' // U+662B <cjk>
	0xEB53: '昰' // U+6630 <cjk>
	0xEB54: '昱' // U+6631 <cjk>
	0xEB55: '昳' // U+6633 <cjk>
	0xEB56: '曻' // U+66FB <cjk>
	0xEB57: '晈' // U+6648 <cjk>
	0xEB58: '晌' // U+664C <cjk>
	0xEB59: '𣇄' // U+231C4 <cjk>
	0xEB5A: '晙' // U+6659 <cjk>
	0xEB5B: '晚' // U+665A <cjk>
	0xEB5C: '晡' // U+6661 <cjk>
	0xEB5D: '晥' // U+6665 <cjk>
	0xEB5E: '晳' // U+6673 <cjk>
	0xEB5F: '晷' // U+6677 <cjk>
	0xEB60: '晸' // U+6678 <cjk>
	0xEB61: '暍' // U+668D <cjk>
	0xEB62: '暑' // U+FA43 CJK COMPATIBILITY IDEOGRAPH-FA43
	0xEB63: '暠' // U+66A0 <cjk>
	0xEB64: '暲' // U+66B2 <cjk>
	0xEB65: '暻' // U+66BB <cjk>
	0xEB66: '曆' // U+66C6 <cjk>
	0xEB67: '曈' // U+66C8 <cjk>
	0xEB68: '㬢' // U+3B22 <cjk>
	0xEB69: '曛' // U+66DB <cjk>
	0xEB6A: '曨' // U+66E8 <cjk>
	0xEB6B: '曺' // U+66FA <cjk>
	0xEB6C: '朓' // U+6713 <cjk>
	0xEB6D: '朗' // U+F929 CJK COMPATIBILITY IDEOGRAPH-F929
	0xEB6E: '朳' // U+6733 <cjk>
	0xEB6F: '杦' // U+6766 <cjk>
	0xEB70: '杇' // U+6747 <cjk>
	0xEB71: '杈' // U+6748 <cjk>
	0xEB72: '杻' // U+677B <cjk>
	0xEB73: '极' // U+6781 <cjk>
	0xEB74: '枓' // U+6793 <cjk>
	0xEB75: '枘' // U+6798 <cjk>
	0xEB76: '枛' // U+679B <cjk>
	0xEB77: '枻' // U+67BB <cjk>
	0xEB78: '柹' // U+67F9 <cjk>
	0xEB79: '柀' // U+67C0 <cjk>
	0xEB7A: '柗' // U+67D7 <cjk>
	0xEB7B: '柼' // U+67FC <cjk>
	0xEB7C: '栁' // U+6801 <cjk>
	0xEB7D: '桒' // U+6852 <cjk>
	0xEB7E: '栝' // U+681D <cjk>
	0xEB80: '栬' // U+682C <cjk>
	0xEB81: '栱' // U+6831 <cjk>
	0xEB82: '桛' // U+685B <cjk>
	0xEB83: '桲' // U+6872 <cjk>
	0xEB84: '桵' // U+6875 <cjk>
	0xEB85: '梅' // U+FA44 CJK COMPATIBILITY IDEOGRAPH-FA44
	0xEB86: '梣' // U+68A3 <cjk>
	0xEB87: '梥' // U+68A5 <cjk>
	0xEB88: '梲' // U+68B2 <cjk>
	0xEB89: '棈' // U+68C8 <cjk>
	0xEB8A: '棐' // U+68D0 <cjk>
	0xEB8B: '棨' // U+68E8 <cjk>
	0xEB8C: '棭' // U+68ED <cjk>
	0xEB8D: '棰' // U+68F0 <cjk>
	0xEB8E: '棱' // U+68F1 <cjk>
	0xEB8F: '棼' // U+68FC <cjk>
	0xEB90: '椊' // U+690A <cjk>
	0xEB91: '楉' // U+6949 <cjk>
	0xEB92: '𣗄' // U+235C4 <cjk>
	0xEB93: '椵' // U+6935 <cjk>
	0xEB94: '楂' // U+6942 <cjk>
	0xEB95: '楗' // U+6957 <cjk>
	0xEB96: '楣' // U+6963 <cjk>
	0xEB97: '楤' // U+6964 <cjk>
	0xEB98: '楨' // U+6968 <cjk>
	0xEB99: '榀' // U+6980 <cjk>
	0xEB9A: '﨔' // U+FA14 CJK COMPATIBILITY IDEOGRAPH-FA14
	0xEB9B: '榥' // U+69A5 <cjk>
	0xEB9C: '榭' // U+69AD <cjk>
	0xEB9D: '槏' // U+69CF <cjk>
	0xEB9E: '㮶' // U+3BB6 <cjk>
	0xEB9F: '㯃' // U+3BC3 <cjk>
	0xEBA0: '槢' // U+69E2 <cjk>
	0xEBA1: '槩' // U+69E9 <cjk>
	0xEBA2: '槪' // U+69EA <cjk>
	0xEBA3: '槵' // U+69F5 <cjk>
	0xEBA4: '槶' // U+69F6 <cjk>
	0xEBA5: '樏' // U+6A0F <cjk>
	0xEBA6: '樕' // U+6A15 <cjk>
	0xEBA7: '𣜿' // U+2373F <cjk>
	0xEBA8: '樻' // U+6A3B <cjk>
	0xEBA9: '樾' // U+6A3E <cjk>
	0xEBAA: '橅' // U+6A45 <cjk>
	0xEBAB: '橐' // U+6A50 <cjk>
	0xEBAC: '橖' // U+6A56 <cjk>
	0xEBAD: '橛' // U+6A5B <cjk>
	0xEBAE: '橫' // U+6A6B <cjk>
	0xEBAF: '橳' // U+6A73 <cjk>
	0xEBB0: '𣝣' // U+23763 <cjk>
	0xEBB1: '檉' // U+6A89 <cjk>
	0xEBB2: '檔' // U+6A94 <cjk>
	0xEBB3: '檝' // U+6A9D <cjk>
	0xEBB4: '檞' // U+6A9E <cjk>
	0xEBB5: '檥' // U+6AA5 <cjk>
	0xEBB6: '櫤' // U+6AE4 <cjk>
	0xEBB7: '櫧' // U+6AE7 <cjk>
	0xEBB8: '㰏' // U+3C0F <cjk>
	0xEBB9: '欄' // U+F91D CJK COMPATIBILITY IDEOGRAPH-F91D
	0xEBBA: '欛' // U+6B1B <cjk>
	0xEBBB: '欞' // U+6B1E <cjk>
	0xEBBC: '欬' // U+6B2C <cjk>
	0xEBBD: '欵' // U+6B35 <cjk>
	0xEBBE: '歆' // U+6B46 <cjk>
	0xEBBF: '歖' // U+6B56 <cjk>
	0xEBC0: '歠' // U+6B60 <cjk>
	0xEBC1: '步' // U+6B65 <cjk>
	0xEBC2: '歧' // U+6B67 <cjk>
	0xEBC3: '歷' // U+6B77 <cjk>
	0xEBC4: '殂' // U+6B82 <cjk>
	0xEBC5: '殩' // U+6BA9 <cjk>
	0xEBC6: '殭' // U+6BAD <cjk>
	0xEBC7: '殺' // U+F970 CJK COMPATIBILITY IDEOGRAPH-F970
	0xEBC8: '每' // U+6BCF <cjk>
	0xEBC9: '毖' // U+6BD6 <cjk>
	0xEBCA: '毗' // U+6BD7 <cjk>
	0xEBCB: '毿' // U+6BFF <cjk>
	0xEBCC: '氅' // U+6C05 <cjk>
	0xEBCD: '氐' // U+6C10 <cjk>
	0xEBCE: '氳' // U+6C33 <cjk>
	0xEBCF: '汙' // U+6C59 <cjk>
	0xEBD0: '汜' // U+6C5C <cjk>
	0xEBD1: '沪' // U+6CAA <cjk>
	0xEBD2: '汴' // U+6C74 <cjk>
	0xEBD3: '汶' // U+6C76 <cjk>
	0xEBD4: '沅' // U+6C85 <cjk>
	0xEBD5: '沆' // U+6C86 <cjk>
	0xEBD6: '沘' // U+6C98 <cjk>
	0xEBD7: '沜' // U+6C9C <cjk>
	0xEBD8: '泻' // U+6CFB <cjk>
	0xEBD9: '泆' // U+6CC6 <cjk>
	0xEBDA: '泔' // U+6CD4 <cjk>
	0xEBDB: '泠' // U+6CE0 <cjk>
	0xEBDC: '泫' // U+6CEB <cjk>
	0xEBDD: '泮' // U+6CEE <cjk>
	0xEBDE: '𣳾' // U+23CFE <cjk>
	0xEBDF: '洄' // U+6D04 <cjk>
	0xEBE0: '洎' // U+6D0E <cjk>
	0xEBE1: '洮' // U+6D2E <cjk>
	0xEBE2: '洱' // U+6D31 <cjk>
	0xEBE3: '洹' // U+6D39 <cjk>
	0xEBE4: '洿' // U+6D3F <cjk>
	0xEBE5: '浘' // U+6D58 <cjk>
	0xEBE6: '浥' // U+6D65 <cjk>
	0xEBE7: '海' // U+FA45 CJK COMPATIBILITY IDEOGRAPH-FA45
	0xEBE8: '涂' // U+6D82 <cjk>
	0xEBE9: '涇' // U+6D87 <cjk>
	0xEBEA: '涉' // U+6D89 <cjk>
	0xEBEB: '涔' // U+6D94 <cjk>
	0xEBEC: '涪' // U+6DAA <cjk>
	0xEBED: '涬' // U+6DAC <cjk>
	0xEBEE: '涿' // U+6DBF <cjk>
	0xEBEF: '淄' // U+6DC4 <cjk>
	0xEBF0: '淖' // U+6DD6 <cjk>
	0xEBF1: '淚' // U+6DDA <cjk>
	0xEBF2: '淛' // U+6DDB <cjk>
	0xEBF3: '淝' // U+6DDD <cjk>
	0xEBF4: '淼' // U+6DFC <cjk>
	0xEBF5: '渚' // U+FA46 CJK COMPATIBILITY IDEOGRAPH-FA46
	0xEBF6: '渴' // U+6E34 <cjk>
	0xEBF7: '湄' // U+6E44 <cjk>
	0xEBF8: '湜' // U+6E5C <cjk>
	0xEBF9: '湞' // U+6E5E <cjk>
	0xEBFA: '溫' // U+6EAB <cjk>
	0xEBFB: '溱' // U+6EB1 <cjk>
	0xEBFC: '滁' // U+6EC1 <cjk>
	0xEC40: '滇' // U+6EC7 <cjk>
	0xEC41: '滎' // U+6ECE <cjk>
	0xEC42: '漐' // U+6F10 <cjk>
	0xEC43: '漚' // U+6F1A <cjk>
	0xEC44: '漢' // U+FA47 CJK COMPATIBILITY IDEOGRAPH-FA47
	0xEC45: '漪' // U+6F2A <cjk>
	0xEC46: '漯' // U+6F2F <cjk>
	0xEC47: '漳' // U+6F33 <cjk>
	0xEC48: '潑' // U+6F51 <cjk>
	0xEC49: '潙' // U+6F59 <cjk>
	0xEC4A: '潞' // U+6F5E <cjk>
	0xEC4B: '潡' // U+6F61 <cjk>
	0xEC4C: '潢' // U+6F62 <cjk>
	0xEC4D: '潾' // U+6F7E <cjk>
	0xEC4E: '澈' // U+6F88 <cjk>
	0xEC4F: '澌' // U+6F8C <cjk>
	0xEC50: '澍' // U+6F8D <cjk>
	0xEC51: '澔' // U+6F94 <cjk>
	0xEC52: '澠' // U+6FA0 <cjk>
	0xEC53: '澧' // U+6FA7 <cjk>
	0xEC54: '澶' // U+6FB6 <cjk>
	0xEC55: '澼' // U+6FBC <cjk>
	0xEC56: '濇' // U+6FC7 <cjk>
	0xEC57: '濊' // U+6FCA <cjk>
	0xEC58: '濹' // U+6FF9 <cjk>
	0xEC59: '濰' // U+6FF0 <cjk>
	0xEC5A: '濵' // U+6FF5 <cjk>
	0xEC5B: '瀅' // U+7005 <cjk>
	0xEC5C: '瀆' // U+7006 <cjk>
	0xEC5D: '瀨' // U+7028 <cjk>
	0xEC5E: '灊' // U+704A <cjk>
	0xEC5F: '灝' // U+705D <cjk>
	0xEC60: '灞' // U+705E <cjk>
	0xEC61: '灎' // U+704E <cjk>
	0xEC62: '灤' // U+7064 <cjk>
	0xEC63: '灵' // U+7075 <cjk>
	0xEC64: '炅' // U+7085 <cjk>
	0xEC65: '炤' // U+70A4 <cjk>
	0xEC66: '炫' // U+70AB <cjk>
	0xEC67: '炷' // U+70B7 <cjk>
	0xEC68: '烔' // U+70D4 <cjk>
	0xEC69: '烘' // U+70D8 <cjk>
	0xEC6A: '烤' // U+70E4 <cjk>
	0xEC6B: '焏' // U+710F <cjk>
	0xEC6C: '焫' // U+712B <cjk>
	0xEC6D: '焞' // U+711E <cjk>
	0xEC6E: '焠' // U+7120 <cjk>
	0xEC6F: '焮' // U+712E <cjk>
	0xEC70: '焰' // U+7130 <cjk>
	0xEC71: '煆' // U+7146 <cjk>
	0xEC72: '煇' // U+7147 <cjk>
	0xEC73: '煑' // U+7151 <cjk>
	0xEC74: '煮' // U+FA48 CJK COMPATIBILITY IDEOGRAPH-FA48
	0xEC75: '煒' // U+7152 <cjk>
	0xEC76: '煜' // U+715C <cjk>
	0xEC77: '煠' // U+7160 <cjk>
	0xEC78: '煨' // U+7168 <cjk>
	0xEC79: '凞' // U+FA15 CJK COMPATIBILITY IDEOGRAPH-FA15
	0xEC7A: '熅' // U+7185 <cjk>
	0xEC7B: '熇' // U+7187 <cjk>
	0xEC7C: '熒' // U+7192 <cjk>
	0xEC7D: '燁' // U+71C1 <cjk>
	0xEC7E: '熺' // U+71BA <cjk>
	0xEC80: '燄' // U+71C4 <cjk>
	0xEC81: '燾' // U+71FE <cjk>
	0xEC82: '爀' // U+7200 <cjk>
	0xEC83: '爕' // U+7215 <cjk>
	0xEC84: '牕' // U+7255 <cjk>
	0xEC85: '牖' // U+7256 <cjk>
	0xEC86: '㸿' // U+3E3F <cjk>
	0xEC87: '犍' // U+728D <cjk>
	0xEC88: '犛' // U+729B <cjk>
	0xEC89: '犾' // U+72BE <cjk>
	0xEC8A: '狀' // U+72C0 <cjk>
	0xEC8B: '狻' // U+72FB <cjk>
	0xEC8C: '𤟱' // U+247F1 <cjk>
	0xEC8D: '猧' // U+7327 <cjk>
	0xEC8E: '猨' // U+7328 <cjk>
	0xEC8F: '猪' // U+FA16 CJK COMPATIBILITY IDEOGRAPH-FA16
	0xEC90: '獐' // U+7350 <cjk>
	0xEC91: '獦' // U+7366 <cjk>
	0xEC92: '獼' // U+737C <cjk>
	0xEC93: '玕' // U+7395 <cjk>
	0xEC94: '玟' // U+739F <cjk>
	0xEC95: '玠' // U+73A0 <cjk>
	0xEC96: '玢' // U+73A2 <cjk>
	0xEC97: '玦' // U+73A6 <cjk>
	0xEC98: '玫' // U+73AB <cjk>
	0xEC99: '珉' // U+73C9 <cjk>
	0xEC9A: '珏' // U+73CF <cjk>
	0xEC9B: '珖' // U+73D6 <cjk>
	0xEC9C: '珙' // U+73D9 <cjk>
	0xEC9D: '珣' // U+73E3 <cjk>
	0xEC9E: '珩' // U+73E9 <cjk>
	0xEC9F: '琇' // U+7407 <cjk>
	0xECA0: '琊' // U+740A <cjk>
	0xECA1: '琚' // U+741A <cjk>
	0xECA2: '琛' // U+741B <cjk>
	0xECA3: '琢' // U+FA4A CJK COMPATIBILITY IDEOGRAPH-FA4A
	0xECA4: '琦' // U+7426 <cjk>
	0xECA5: '琨' // U+7428 <cjk>
	0xECA6: '琪' // U+742A <cjk>
	0xECA7: '琫' // U+742B <cjk>
	0xECA8: '琬' // U+742C <cjk>
	0xECA9: '琮' // U+742E <cjk>
	0xECAA: '琯' // U+742F <cjk>
	0xECAB: '琰' // U+7430 <cjk>
	0xECAC: '瑄' // U+7444 <cjk>
	0xECAD: '瑆' // U+7446 <cjk>
	0xECAE: '瑇' // U+7447 <cjk>
	0xECAF: '瑋' // U+744B <cjk>
	0xECB0: '瑗' // U+7457 <cjk>
	0xECB1: '瑢' // U+7462 <cjk>
	0xECB2: '瑫' // U+746B <cjk>
	0xECB3: '瑭' // U+746D <cjk>
	0xECB4: '璆' // U+7486 <cjk>
	0xECB5: '璇' // U+7487 <cjk>
	0xECB6: '璉' // U+7489 <cjk>
	0xECB7: '璘' // U+7498 <cjk>
	0xECB8: '璜' // U+749C <cjk>
	0xECB9: '璟' // U+749F <cjk>
	0xECBA: '璣' // U+74A3 <cjk>
	0xECBB: '璐' // U+7490 <cjk>
	0xECBC: '璦' // U+74A6 <cjk>
	0xECBD: '璨' // U+74A8 <cjk>
	0xECBE: '璩' // U+74A9 <cjk>
	0xECBF: '璵' // U+74B5 <cjk>
	0xECC0: '璿' // U+74BF <cjk>
	0xECC1: '瓈' // U+74C8 <cjk>
	0xECC2: '瓉' // U+74C9 <cjk>
	0xECC3: '瓚' // U+74DA <cjk>
	0xECC4: '瓿' // U+74FF <cjk>
	0xECC5: '甁' // U+7501 <cjk>
	0xECC6: '甗' // U+7517 <cjk>
	0xECC7: '甯' // U+752F <cjk>
	0xECC8: '畯' // U+756F <cjk>
	0xECC9: '畹' // U+7579 <cjk>
	0xECCA: '疒' // U+7592 <cjk>
	0xECCB: '㽲' // U+3F72 <cjk>
	0xECCC: '痎' // U+75CE <cjk>
	0xECCD: '痤' // U+75E4 <cjk>
	0xECCE: '瘀' // U+7600 <cjk>
	0xECCF: '瘂' // U+7602 <cjk>
	0xECD0: '瘈' // U+7608 <cjk>
	0xECD1: '瘕' // U+7615 <cjk>
	0xECD2: '瘖' // U+7616 <cjk>
	0xECD3: '瘙' // U+7619 <cjk>
	0xECD4: '瘞' // U+761E <cjk>
	0xECD5: '瘭' // U+762D <cjk>
	0xECD6: '瘵' // U+7635 <cjk>
	0xECD7: '癃' // U+7643 <cjk>
	0xECD8: '癋' // U+764B <cjk>
	0xECD9: '癤' // U+7664 <cjk>
	0xECDA: '癥' // U+7665 <cjk>
	0xECDB: '癭' // U+766D <cjk>
	0xECDC: '癯' // U+766F <cjk>
	0xECDD: '癱' // U+7671 <cjk>
	0xECDE: '皁' // U+7681 <cjk>
	0xECDF: '皛' // U+769B <cjk>
	0xECE0: '皝' // U+769D <cjk>
	0xECE1: '皞' // U+769E <cjk>
	0xECE2: '皦' // U+76A6 <cjk>
	0xECE3: '皪' // U+76AA <cjk>
	0xECE4: '皶' // U+76B6 <cjk>
	0xECE5: '盅' // U+76C5 <cjk>
	0xECE6: '盌' // U+76CC <cjk>
	0xECE7: '盎' // U+76CE <cjk>
	0xECE8: '盔' // U+76D4 <cjk>
	0xECE9: '盦' // U+76E6 <cjk>
	0xECEA: '盱' // U+76F1 <cjk>
	0xECEB: '盼' // U+76FC <cjk>
	0xECEC: '眊' // U+770A <cjk>
	0xECED: '眙' // U+7719 <cjk>
	0xECEE: '眴' // U+7734 <cjk>
	0xECEF: '眶' // U+7736 <cjk>
	0xECF0: '睆' // U+7746 <cjk>
	0xECF1: '睍' // U+774D <cjk>
	0xECF2: '睎' // U+774E <cjk>
	0xECF3: '睜' // U+775C <cjk>
	0xECF4: '睟' // U+775F <cjk>
	0xECF5: '睢' // U+7762 <cjk>
	0xECF6: '睺' // U+777A <cjk>
	0xECF7: '瞀' // U+7780 <cjk>
	0xECF8: '瞔' // U+7794 <cjk>
	0xECF9: '瞪' // U+77AA <cjk>
	0xECFA: '矠' // U+77E0 <cjk>
	0xECFB: '砭' // U+782D <cjk>
	0xECFC: '𥒎' // U+2548E <cjk>
	0xED40: '硃' // U+7843 <cjk>
	0xED41: '硎' // U+784E <cjk>
	0xED42: '硏' // U+784F <cjk>
	0xED43: '硑' // U+7851 <cjk>
	0xED44: '硨' // U+7868 <cjk>
	0xED45: '确' // U+786E <cjk>
	0xED46: '碑' // U+FA4B CJK COMPATIBILITY IDEOGRAPH-FA4B
	0xED47: '碰' // U+78B0 <cjk>
	0xED48: '𥔎' // U+2550E <cjk>
	0xED49: '碭' // U+78AD <cjk>
	0xED4A: '磤' // U+78E4 <cjk>
	0xED4B: '磲' // U+78F2 <cjk>
	0xED4C: '礀' // U+7900 <cjk>
	0xED4D: '磷' // U+78F7 <cjk>
	0xED4E: '礜' // U+791C <cjk>
	0xED4F: '礮' // U+792E <cjk>
	0xED50: '礱' // U+7931 <cjk>
	0xED51: '礴' // U+7934 <cjk>
	0xED52: '社' // U+FA4C CJK COMPATIBILITY IDEOGRAPH-FA4C
	0xED53: '祉' // U+FA4D CJK COMPATIBILITY IDEOGRAPH-FA4D
	0xED54: '祅' // U+7945 <cjk>
	0xED55: '祆' // U+7946 <cjk>
	0xED56: '祈' // U+FA4E CJK COMPATIBILITY IDEOGRAPH-FA4E
	0xED57: '祐' // U+FA4F CJK COMPATIBILITY IDEOGRAPH-FA4F
	0xED58: '祖' // U+FA50 CJK COMPATIBILITY IDEOGRAPH-FA50
	0xED59: '祜' // U+795C <cjk>
	0xED5A: '祝' // U+FA51 CJK COMPATIBILITY IDEOGRAPH-FA51
	0xED5B: '神' // U+FA19 CJK COMPATIBILITY IDEOGRAPH-FA19
	0xED5C: '祥' // U+FA1A CJK COMPATIBILITY IDEOGRAPH-FA1A
	0xED5D: '祹' // U+7979 <cjk>
	0xED5E: '禍' // U+FA52 CJK COMPATIBILITY IDEOGRAPH-FA52
	0xED5F: '禎' // U+FA53 CJK COMPATIBILITY IDEOGRAPH-FA53
	0xED60: '福' // U+FA1B CJK COMPATIBILITY IDEOGRAPH-FA1B
	0xED61: '禘' // U+7998 <cjk>
	0xED62: '禱' // U+79B1 <cjk>
	0xED63: '禸' // U+79B8 <cjk>
	0xED64: '秈' // U+79C8 <cjk>
	0xED65: '秊' // U+79CA <cjk>
	0xED66: '𥝱' // U+25771 <cjk>
	0xED67: '秔' // U+79D4 <cjk>
	0xED68: '秞' // U+79DE <cjk>
	0xED69: '秫' // U+79EB <cjk>
	0xED6A: '秭' // U+79ED <cjk>
	0xED6B: '稃' // U+7A03 <cjk>
	0xED6C: '穀' // U+FA54 CJK COMPATIBILITY IDEOGRAPH-FA54
	0xED6D: '稹' // U+7A39 <cjk>
	0xED6E: '穝' // U+7A5D <cjk>
	0xED6F: '穭' // U+7A6D <cjk>
	0xED70: '突' // U+FA55 CJK COMPATIBILITY IDEOGRAPH-FA55
	0xED71: '窅' // U+7A85 <cjk>
	0xED72: '窠' // U+7AA0 <cjk>
	0xED73: '𥧄' // U+259C4 <cjk>
	0xED74: '窳' // U+7AB3 <cjk>
	0xED75: '窻' // U+7ABB <cjk>
	0xED76: '竎' // U+7ACE <cjk>
	0xED77: '竫' // U+7AEB <cjk>
	0xED78: '竽' // U+7AFD <cjk>
	0xED79: '笒' // U+7B12 <cjk>
	0xED7A: '笭' // U+7B2D <cjk>
	0xED7B: '笻' // U+7B3B <cjk>
	0xED7C: '筇' // U+7B47 <cjk>
	0xED7D: '筎' // U+7B4E <cjk>
	0xED7E: '筠' // U+7B60 <cjk>
	0xED80: '筭' // U+7B6D <cjk>
	0xED81: '筯' // U+7B6F <cjk>
	0xED82: '筲' // U+7B72 <cjk>
	0xED83: '箞' // U+7B9E <cjk>
	0xED84: '節' // U+FA56 CJK COMPATIBILITY IDEOGRAPH-FA56
	0xED85: '篗' // U+7BD7 <cjk>
	0xED86: '篙' // U+7BD9 <cjk>
	0xED87: '簁' // U+7C01 <cjk>
	0xED88: '簱' // U+7C31 <cjk>
	0xED89: '簞' // U+7C1E <cjk>
	0xED8A: '簠' // U+7C20 <cjk>
	0xED8B: '簳' // U+7C33 <cjk>
	0xED8C: '簶' // U+7C36 <cjk>
	0xED8D: '䉤' // U+4264 <cjk>
	0xED8E: '𥶡' // U+25DA1 <cjk>
	0xED8F: '籙' // U+7C59 <cjk>
	0xED90: '籭' // U+7C6D <cjk>
	0xED91: '籹' // U+7C79 <cjk>
	0xED92: '粏' // U+7C8F <cjk>
	0xED93: '粔' // U+7C94 <cjk>
	0xED94: '粠' // U+7CA0 <cjk>
	0xED95: '粼' // U+7CBC <cjk>
	0xED96: '糕' // U+7CD5 <cjk>
	0xED97: '糙' // U+7CD9 <cjk>
	0xED98: '糝' // U+7CDD <cjk>
	0xED99: '紇' // U+7D07 <cjk>
	0xED9A: '紈' // U+7D08 <cjk>
	0xED9B: '紓' // U+7D13 <cjk>
	0xED9C: '紝' // U+7D1D <cjk>
	0xED9D: '紣' // U+7D23 <cjk>
	0xED9E: '紱' // U+7D31 <cjk>
	0xED9F: '絁' // U+7D41 <cjk>
	0xEDA0: '絈' // U+7D48 <cjk>
	0xEDA1: '絓' // U+7D53 <cjk>
	0xEDA2: '絜' // U+7D5C <cjk>
	0xEDA3: '絺' // U+7D7A <cjk>
	0xEDA4: '綃' // U+7D83 <cjk>
	0xEDA5: '綋' // U+7D8B <cjk>
	0xEDA6: '綠' // U+7DA0 <cjk>
	0xEDA7: '綦' // U+7DA6 <cjk>
	0xEDA8: '緂' // U+7DC2 <cjk>
	0xEDA9: '緌' // U+7DCC <cjk>
	0xEDAA: '緖' // U+7DD6 <cjk>
	0xEDAB: '緣' // U+7DE3 <cjk>
	0xEDAC: '練' // U+FA57 CJK COMPATIBILITY IDEOGRAPH-FA57
	0xEDAD: '縨' // U+7E28 <cjk>
	0xEDAE: '縈' // U+7E08 <cjk>
	0xEDAF: '縑' // U+7E11 <cjk>
	0xEDB0: '縕' // U+7E15 <cjk>
	0xEDB1: '繁' // U+FA59 CJK COMPATIBILITY IDEOGRAPH-FA59
	0xEDB2: '繇' // U+7E47 <cjk>
	0xEDB3: '繒' // U+7E52 <cjk>
	0xEDB4: '繡' // U+7E61 <cjk>
	0xEDB5: '纊' // U+7E8A <cjk>
	0xEDB6: '纍' // U+7E8D <cjk>
	0xEDB7: '罇' // U+7F47 <cjk>
	0xEDB8: '署' // U+FA5A CJK COMPATIBILITY IDEOGRAPH-FA5A
	0xEDB9: '羑' // U+7F91 <cjk>
	0xEDBA: '羗' // U+7F97 <cjk>
	0xEDBB: '羿' // U+7FBF <cjk>
	0xEDBC: '翎' // U+7FCE <cjk>
	0xEDBD: '翛' // U+7FDB <cjk>
	0xEDBE: '翟' // U+7FDF <cjk>
	0xEDBF: '翬' // U+7FEC <cjk>
	0xEDC0: '翮' // U+7FEE <cjk>
	0xEDC1: '翺' // U+7FFA <cjk>
	0xEDC2: '者' // U+FA5B CJK COMPATIBILITY IDEOGRAPH-FA5B
	0xEDC3: '耔' // U+8014 <cjk>
	0xEDC4: '耦' // U+8026 <cjk>
	0xEDC5: '耵' // U+8035 <cjk>
	0xEDC6: '耷' // U+8037 <cjk>
	0xEDC7: '耼' // U+803C <cjk>
	0xEDC8: '胊' // U+80CA <cjk>
	0xEDC9: '胗' // U+80D7 <cjk>
	0xEDCA: '胠' // U+80E0 <cjk>
	0xEDCB: '胳' // U+80F3 <cjk>
	0xEDCC: '脘' // U+8118 <cjk>
	0xEDCD: '腊' // U+814A <cjk>
	0xEDCE: '腠' // U+8160 <cjk>
	0xEDCF: '腧' // U+8167 <cjk>
	0xEDD0: '腨' // U+8168 <cjk>
	0xEDD1: '腭' // U+816D <cjk>
	0xEDD2: '膻' // U+81BB <cjk>
	0xEDD3: '臊' // U+81CA <cjk>
	0xEDD4: '臏' // U+81CF <cjk>
	0xEDD5: '臗' // U+81D7 <cjk>
	0xEDD6: '臭' // U+FA5C CJK COMPATIBILITY IDEOGRAPH-FA5C
	0xEDD7: '䑓' // U+4453 <cjk>
	0xEDD8: '䑛' // U+445B <cjk>
	0xEDD9: '艠' // U+8260 <cjk>
	0xEDDA: '艴' // U+8274 <cjk>
	0xEDDB: '𦫿' // U+26AFF <cjk>
	0xEDDC: '芎' // U+828E <cjk>
	0xEDDD: '芡' // U+82A1 <cjk>
	0xEDDE: '芣' // U+82A3 <cjk>
	0xEDDF: '芤' // U+82A4 <cjk>
	0xEDE0: '芩' // U+82A9 <cjk>
	0xEDE1: '芮' // U+82AE <cjk>
	0xEDE2: '芷' // U+82B7 <cjk>
	0xEDE3: '芾' // U+82BE <cjk>
	0xEDE4: '芿' // U+82BF <cjk>
	0xEDE5: '苆' // U+82C6 <cjk>
	0xEDE6: '苕' // U+82D5 <cjk>
	0xEDE7: '苽' // U+82FD <cjk>
	0xEDE8: '苾' // U+82FE <cjk>
	0xEDE9: '茀' // U+8300 <cjk>
	0xEDEA: '茁' // U+8301 <cjk>
	0xEDEB: '荢' // U+8362 <cjk>
	0xEDEC: '茢' // U+8322 <cjk>
	0xEDED: '茭' // U+832D <cjk>
	0xEDEE: '茺' // U+833A <cjk>
	0xEDEF: '荃' // U+8343 <cjk>
	0xEDF0: '荇' // U+8347 <cjk>
	0xEDF1: '荑' // U+8351 <cjk>
	0xEDF2: '荕' // U+8355 <cjk>
	0xEDF3: '荽' // U+837D <cjk>
	0xEDF4: '莆' // U+8386 <cjk>
	0xEDF5: '莒' // U+8392 <cjk>
	0xEDF6: '莘' // U+8398 <cjk>
	0xEDF7: '莧' // U+83A7 <cjk>
	0xEDF8: '莩' // U+83A9 <cjk>
	0xEDF9: '莿' // U+83BF <cjk>
	0xEDFA: '菀' // U+83C0 <cjk>
	0xEDFB: '菇' // U+83C7 <cjk>
	0xEDFC: '菏' // U+83CF <cjk>
	0xEE40: '菑' // U+83D1 <cjk>
	0xEE41: '菡' // U+83E1 <cjk>
	0xEE42: '菪' // U+83EA <cjk>
	0xEE43: '萁' // U+8401 <cjk>
	0xEE44: '萆' // U+8406 <cjk>
	0xEE45: '萊' // U+840A <cjk>
	0xEE46: '著' // U+FA5F CJK COMPATIBILITY IDEOGRAPH-FA5F
	0xEE47: '葈' // U+8448 <cjk>
	0xEE48: '葟' // U+845F <cjk>
	0xEE49: '葰' // U+8470 <cjk>
	0xEE4A: '葳' // U+8473 <cjk>
	0xEE4B: '蒅' // U+8485 <cjk>
	0xEE4C: '蒞' // U+849E <cjk>
	0xEE4D: '蒯' // U+84AF <cjk>
	0xEE4E: '蒴' // U+84B4 <cjk>
	0xEE4F: '蒺' // U+84BA <cjk>
	0xEE50: '蓀' // U+84C0 <cjk>
	0xEE51: '蓂' // U+84C2 <cjk>
	0xEE52: '𦹀' // U+26E40 <cjk>
	0xEE53: '蔲' // U+8532 <cjk>
	0xEE54: '蔞' // U+851E <cjk>
	0xEE55: '蔣' // U+8523 <cjk>
	0xEE56: '蔯' // U+852F <cjk>
	0xEE57: '蕙' // U+8559 <cjk>
	0xEE58: '蕤' // U+8564 <cjk>
	0xEE59: '﨟' // U+FA1F CJK COMPATIBILITY IDEOGRAPH-FA1F
	0xEE5A: '薭' // U+85AD <cjk>
	0xEE5B: '蕺' // U+857A <cjk>
	0xEE5C: '薌' // U+858C <cjk>
	0xEE5D: '薏' // U+858F <cjk>
	0xEE5E: '薢' // U+85A2 <cjk>
	0xEE5F: '薰' // U+85B0 <cjk>
	0xEE60: '藋' // U+85CB <cjk>
	0xEE61: '藎' // U+85CE <cjk>
	0xEE62: '藭' // U+85ED <cjk>
	0xEE63: '蘒' // U+8612 <cjk>
	0xEE64: '藿' // U+85FF <cjk>
	0xEE65: '蘄' // U+8604 <cjk>
	0xEE66: '蘅' // U+8605 <cjk>
	0xEE67: '蘐' // U+8610 <cjk>
	0xEE68: '𧃴' // U+270F4 <cjk>
	0xEE69: '蘘' // U+8618 <cjk>
	0xEE6A: '蘩' // U+8629 <cjk>
	0xEE6B: '蘸' // U+8638 <cjk>
	0xEE6C: '虗' // U+8657 <cjk>
	0xEE6D: '虛' // U+865B <cjk>
	0xEE6E: '虜' // U+F936 CJK COMPATIBILITY IDEOGRAPH-F936
	0xEE6F: '虢' // U+8662 <cjk>
	0xEE70: '䖝' // U+459D <cjk>
	0xEE71: '虬' // U+866C <cjk>
	0xEE72: '虵' // U+8675 <cjk>
	0xEE73: '蚘' // U+8698 <cjk>
	0xEE74: '蚸' // U+86B8 <cjk>
	0xEE75: '蛺' // U+86FA <cjk>
	0xEE76: '蛼' // U+86FC <cjk>
	0xEE77: '蛽' // U+86FD <cjk>
	0xEE78: '蜋' // U+870B <cjk>
	0xEE79: '蝱' // U+8771 <cjk>
	0xEE7A: '螇' // U+8787 <cjk>
	0xEE7B: '螈' // U+8788 <cjk>
	0xEE7C: '螬' // U+87AC <cjk>
	0xEE7D: '螭' // U+87AD <cjk>
	0xEE7E: '螵' // U+87B5 <cjk>
	0xEE80: '䗪' // U+45EA <cjk>
	0xEE81: '蟖' // U+87D6 <cjk>
	0xEE82: '蟬' // U+87EC <cjk>
	0xEE83: '蠆' // U+8806 <cjk>
	0xEE84: '蠊' // U+880A <cjk>
	0xEE85: '蠐' // U+8810 <cjk>
	0xEE86: '蠔' // U+8814 <cjk>
	0xEE87: '蠟' // U+881F <cjk>
	0xEE88: '袘' // U+8898 <cjk>
	0xEE89: '袪' // U+88AA <cjk>
	0xEE8A: '裊' // U+88CA <cjk>
	0xEE8B: '裎' // U+88CE <cjk>
	0xEE8C: '𧚄' // U+27684 <cjk>
	0xEE8D: '裵' // U+88F5 <cjk>
	0xEE8E: '褜' // U+891C <cjk>
	0xEE8F: '褐' // U+FA60 CJK COMPATIBILITY IDEOGRAPH-FA60
	0xEE90: '褘' // U+8918 <cjk>
	0xEE91: '褙' // U+8919 <cjk>
	0xEE92: '褚' // U+891A <cjk>
	0xEE93: '褧' // U+8927 <cjk>
	0xEE94: '褰' // U+8930 <cjk>
	0xEE95: '褲' // U+8932 <cjk>
	0xEE96: '褹' // U+8939 <cjk>
	0xEE97: '襀' // U+8940 <cjk>
	0xEE98: '覔' // U+8994 <cjk>
	0xEE99: '視' // U+FA61 CJK COMPATIBILITY IDEOGRAPH-FA61
	0xEE9A: '觔' // U+89D4 <cjk>
	0xEE9B: '觥' // U+89E5 <cjk>
	0xEE9C: '觶' // U+89F6 <cjk>
	0xEE9D: '訒' // U+8A12 <cjk>
	0xEE9E: '訕' // U+8A15 <cjk>
	0xEE9F: '訢' // U+8A22 <cjk>
	0xEEA0: '訷' // U+8A37 <cjk>
	0xEEA1: '詇' // U+8A47 <cjk>
	0xEEA2: '詎' // U+8A4E <cjk>
	0xEEA3: '詝' // U+8A5D <cjk>
	0xEEA4: '詡' // U+8A61 <cjk>
	0xEEA5: '詵' // U+8A75 <cjk>
	0xEEA6: '詹' // U+8A79 <cjk>
	0xEEA7: '誧' // U+8AA7 <cjk>
	0xEEA8: '諐' // U+8AD0 <cjk>
	0xEEA9: '諟' // U+8ADF <cjk>
	0xEEAA: '諴' // U+8AF4 <cjk>
	0xEEAB: '諶' // U+8AF6 <cjk>
	0xEEAC: '諸' // U+FA22 CJK COMPATIBILITY IDEOGRAPH-FA22
	0xEEAD: '謁' // U+FA62 CJK COMPATIBILITY IDEOGRAPH-FA62
	0xEEAE: '謹' // U+FA63 CJK COMPATIBILITY IDEOGRAPH-FA63
	0xEEAF: '譆' // U+8B46 <cjk>
	0xEEB0: '譔' // U+8B54 <cjk>
	0xEEB1: '譙' // U+8B59 <cjk>
	0xEEB2: '譩' // U+8B69 <cjk>
	0xEEB3: '讝' // U+8B9D <cjk>
	0xEEB4: '豉' // U+8C49 <cjk>
	0xEEB5: '豨' // U+8C68 <cjk>
	0xEEB6: '賓' // U+FA64 CJK COMPATIBILITY IDEOGRAPH-FA64
	0xEEB7: '賡' // U+8CE1 <cjk>
	0xEEB8: '賴' // U+8CF4 <cjk>
	0xEEB9: '賸' // U+8CF8 <cjk>
	0xEEBA: '賾' // U+8CFE <cjk>
	0xEEBB: '贈' // U+FA65 CJK COMPATIBILITY IDEOGRAPH-FA65
	0xEEBC: '贒' // U+8D12 <cjk>
	0xEEBD: '贛' // U+8D1B <cjk>
	0xEEBE: '趯' // U+8DAF <cjk>
	0xEEBF: '跎' // U+8DCE <cjk>
	0xEEC0: '跑' // U+8DD1 <cjk>
	0xEEC1: '跗' // U+8DD7 <cjk>
	0xEEC2: '踠' // U+8E20 <cjk>
	0xEEC3: '踣' // U+8E23 <cjk>
	0xEEC4: '踽' // U+8E3D <cjk>
	0xEEC5: '蹰' // U+8E70 <cjk>
	0xEEC6: '蹻' // U+8E7B <cjk>
	0xEEC7: '𨉷' // U+28277 <cjk>
	0xEEC8: '軀' // U+8EC0 <cjk>
	0xEEC9: '䡄' // U+4844 <cjk>
	0xEECA: '軺' // U+8EFA <cjk>
	0xEECB: '輞' // U+8F1E <cjk>
	0xEECC: '輭' // U+8F2D <cjk>
	0xEECD: '輶' // U+8F36 <cjk>
	0xEECE: '轔' // U+8F54 <cjk>
	0xEECF: '𨏍' // U+283CD <cjk>
	0xEED0: '辦' // U+8FA6 <cjk>
	0xEED1: '辵' // U+8FB5 <cjk>
	0xEED2: '迤' // U+8FE4 <cjk>
	0xEED3: '迨' // U+8FE8 <cjk>
	0xEED4: '迮' // U+8FEE <cjk>
	0xEED5: '逈' // U+9008 <cjk>
	0xEED6: '逭' // U+902D <cjk>
	0xEED7: '逸' // U+FA67 CJK COMPATIBILITY IDEOGRAPH-FA67
	0xEED8: '邈' // U+9088 <cjk>
	0xEED9: '邕' // U+9095 <cjk>
	0xEEDA: '邗' // U+9097 <cjk>
	0xEEDB: '邙' // U+9099 <cjk>
	0xEEDC: '邛' // U+909B <cjk>
	0xEEDD: '邢' // U+90A2 <cjk>
	0xEEDE: '邳' // U+90B3 <cjk>
	0xEEDF: '邾' // U+90BE <cjk>
	0xEEE0: '郄' // U+90C4 <cjk>
	0xEEE1: '郅' // U+90C5 <cjk>
	0xEEE2: '郇' // U+90C7 <cjk>
	0xEEE3: '郗' // U+90D7 <cjk>
	0xEEE4: '郝' // U+90DD <cjk>
	0xEEE5: '郞' // U+90DE <cjk>
	0xEEE6: '郯' // U+90EF <cjk>
	0xEEE7: '郴' // U+90F4 <cjk>
	0xEEE8: '都' // U+FA26 CJK COMPATIBILITY IDEOGRAPH-FA26
	0xEEE9: '鄔' // U+9114 <cjk>
	0xEEEA: '鄕' // U+9115 <cjk>
	0xEEEB: '鄖' // U+9116 <cjk>
	0xEEEC: '鄢' // U+9122 <cjk>
	0xEEED: '鄣' // U+9123 <cjk>
	0xEEEE: '鄧' // U+9127 <cjk>
	0xEEEF: '鄯' // U+912F <cjk>
	0xEEF0: '鄱' // U+9131 <cjk>
	0xEEF1: '鄴' // U+9134 <cjk>
	0xEEF2: '鄽' // U+913D <cjk>
	0xEEF3: '酈' // U+9148 <cjk>
	0xEEF4: '酛' // U+915B <cjk>
	0xEEF5: '醃' // U+9183 <cjk>
	0xEEF6: '醞' // U+919E <cjk>
	0xEEF7: '醬' // U+91AC <cjk>
	0xEEF8: '醱' // U+91B1 <cjk>
	0xEEF9: '醼' // U+91BC <cjk>
	0xEEFA: '釗' // U+91D7 <cjk>
	0xEEFB: '釻' // U+91FB <cjk>
	0xEEFC: '釤' // U+91E4 <cjk>
	0xEF40: '釥' // U+91E5 <cjk>
	0xEF41: '釭' // U+91ED <cjk>
	0xEF42: '釱' // U+91F1 <cjk>
	0xEF43: '鈇' // U+9207 <cjk>
	0xEF44: '鈐' // U+9210 <cjk>
	0xEF45: '鈸' // U+9238 <cjk>
	0xEF46: '鈹' // U+9239 <cjk>
	0xEF47: '鈺' // U+923A <cjk>
	0xEF48: '鈼' // U+923C <cjk>
	0xEF49: '鉀' // U+9240 <cjk>
	0xEF4A: '鉃' // U+9243 <cjk>
	0xEF4B: '鉏' // U+924F <cjk>
	0xEF4C: '鉸' // U+9278 <cjk>
	0xEF4D: '銈' // U+9288 <cjk>
	0xEF4E: '鋂' // U+92C2 <cjk>
	0xEF4F: '鋋' // U+92CB <cjk>
	0xEF50: '鋌' // U+92CC <cjk>
	0xEF51: '鋓' // U+92D3 <cjk>
	0xEF52: '鋠' // U+92E0 <cjk>
	0xEF53: '鋿' // U+92FF <cjk>
	0xEF54: '錄' // U+9304 <cjk>
	0xEF55: '錟' // U+931F <cjk>
	0xEF56: '錡' // U+9321 <cjk>
	0xEF57: '錥' // U+9325 <cjk>
	0xEF58: '鍈' // U+9348 <cjk>
	0xEF59: '鍉' // U+9349 <cjk>
	0xEF5A: '鍊' // U+934A <cjk>
	0xEF5B: '鍤' // U+9364 <cjk>
	0xEF5C: '鍥' // U+9365 <cjk>
	0xEF5D: '鍪' // U+936A <cjk>
	0xEF5E: '鍰' // U+9370 <cjk>
	0xEF5F: '鎛' // U+939B <cjk>
	0xEF60: '鎣' // U+93A3 <cjk>
	0xEF61: '鎺' // U+93BA <cjk>
	0xEF62: '鏆' // U+93C6 <cjk>
	0xEF63: '鏞' // U+93DE <cjk>
	0xEF64: '鏟' // U+93DF <cjk>
	0xEF65: '鐄' // U+9404 <cjk>
	0xEF66: '鏽' // U+93FD <cjk>
	0xEF67: '鐳' // U+9433 <cjk>
	0xEF68: '鑊' // U+944A <cjk>
	0xEF69: '鑣' // U+9463 <cjk>
	0xEF6A: '鑫' // U+946B <cjk>
	0xEF6B: '鑱' // U+9471 <cjk>
	0xEF6C: '鑲' // U+9472 <cjk>
	0xEF6D: '閎' // U+958E <cjk>
	0xEF6E: '閟' // U+959F <cjk>
	0xEF6F: '閦' // U+95A6 <cjk>
	0xEF70: '閩' // U+95A9 <cjk>
	0xEF71: '閬' // U+95AC <cjk>
	0xEF72: '閶' // U+95B6 <cjk>
	0xEF73: '閽' // U+95BD <cjk>
	0xEF74: '闋' // U+95CB <cjk>
	0xEF75: '闐' // U+95D0 <cjk>
	0xEF76: '闓' // U+95D3 <cjk>
	0xEF77: '䦰' // U+49B0 <cjk>
	0xEF78: '闚' // U+95DA <cjk>
	0xEF79: '闞' // U+95DE <cjk>
	0xEF7A: '陘' // U+9658 <cjk>
	0xEF7B: '隄' // U+9684 <cjk>
	0xEF7C: '隆' // U+F9DC CJK COMPATIBILITY IDEOGRAPH-F9DC
	0xEF7D: '隝' // U+969D <cjk>
	0xEF7E: '隤' // U+96A4 <cjk>
	0xEF80: '隥' // U+96A5 <cjk>
	0xEF81: '雒' // U+96D2 <cjk>
	0xEF82: '雞' // U+96DE <cjk>
	0xEF83: '難' // U+FA68 CJK COMPATIBILITY IDEOGRAPH-FA68
	0xEF84: '雩' // U+96E9 <cjk>
	0xEF85: '雯' // U+96EF <cjk>
	0xEF86: '霳' // U+9733 <cjk>
	0xEF87: '霻' // U+973B <cjk>
	0xEF88: '靍' // U+974D <cjk>
	0xEF89: '靎' // U+974E <cjk>
	0xEF8A: '靏' // U+974F <cjk>
	0xEF8B: '靚' // U+975A <cjk>
	0xEF8C: '靮' // U+976E <cjk>
	0xEF8D: '靳' // U+9773 <cjk>
	0xEF8E: '鞕' // U+9795 <cjk>
	0xEF8F: '鞮' // U+97AE <cjk>
	0xEF90: '鞺' // U+97BA <cjk>
	0xEF91: '韁' // U+97C1 <cjk>
	0xEF92: '韉' // U+97C9 <cjk>
	0xEF93: '韞' // U+97DE <cjk>
	0xEF94: '韛' // U+97DB <cjk>
	0xEF95: '韴' // U+97F4 <cjk>
	0xEF96: '響' // U+FA69 CJK COMPATIBILITY IDEOGRAPH-FA69
	0xEF97: '頊' // U+980A <cjk>
	0xEF98: '頞' // U+981E <cjk>
	0xEF99: '頫' // U+982B <cjk>
	0xEF9A: '頰' // U+9830 <cjk>
	0xEF9B: '頻' // U+FA6A CJK COMPATIBILITY IDEOGRAPH-FA6A
	0xEF9C: '顒' // U+9852 <cjk>
	0xEF9D: '顓' // U+9853 <cjk>
	0xEF9E: '顖' // U+9856 <cjk>
	0xEF9F: '顗' // U+9857 <cjk>
	0xEFA0: '顙' // U+9859 <cjk>
	0xEFA1: '顚' // U+985A <cjk>
	0xEFA2: '類' // U+F9D0 CJK COMPATIBILITY IDEOGRAPH-F9D0
	0xEFA3: '顥' // U+9865 <cjk>
	0xEFA4: '顬' // U+986C <cjk>
	0xEFA5: '颺' // U+98BA <cjk>
	0xEFA6: '飈' // U+98C8 <cjk>
	0xEFA7: '飧' // U+98E7 <cjk>
	0xEFA8: '饘' // U+9958 <cjk>
	0xEFA9: '馞' // U+999E <cjk>
	0xEFAA: '騂' // U+9A02 <cjk>
	0xEFAB: '騃' // U+9A03 <cjk>
	0xEFAC: '騤' // U+9A24 <cjk>
	0xEFAD: '騭' // U+9A2D <cjk>
	0xEFAE: '騮' // U+9A2E <cjk>
	0xEFAF: '騸' // U+9A38 <cjk>
	0xEFB0: '驊' // U+9A4A <cjk>
	0xEFB1: '驎' // U+9A4E <cjk>
	0xEFB2: '驒' // U+9A52 <cjk>
	0xEFB3: '骶' // U+9AB6 <cjk>
	0xEFB4: '髁' // U+9AC1 <cjk>
	0xEFB5: '髃' // U+9AC3 <cjk>
	0xEFB6: '髎' // U+9ACE <cjk>
	0xEFB7: '髖' // U+9AD6 <cjk>
	0xEFB8: '髹' // U+9AF9 <cjk>
	0xEFB9: '鬂' // U+9B02 <cjk>
	0xEFBA: '鬈' // U+9B08 <cjk>
	0xEFBB: '鬠' // U+9B20 <cjk>
	0xEFBC: '䰗' // U+4C17 <cjk>
	0xEFBD: '鬭' // U+9B2D <cjk>
	0xEFBE: '魞' // U+9B5E <cjk>
	0xEFBF: '魹' // U+9B79 <cjk>
	0xEFC0: '魦' // U+9B66 <cjk>
	0xEFC1: '魲' // U+9B72 <cjk>
	0xEFC2: '魵' // U+9B75 <cjk>
	0xEFC3: '鮄' // U+9B84 <cjk>
	0xEFC4: '鮊' // U+9B8A <cjk>
	0xEFC5: '鮏' // U+9B8F <cjk>
	0xEFC6: '鮞' // U+9B9E <cjk>
	0xEFC7: '鮧' // U+9BA7 <cjk>
	0xEFC8: '鯁' // U+9BC1 <cjk>
	0xEFC9: '鯎' // U+9BCE <cjk>
	0xEFCA: '鯥' // U+9BE5 <cjk>
	0xEFCB: '鯸' // U+9BF8 <cjk>
	0xEFCC: '鯽' // U+9BFD <cjk>
	0xEFCD: '鰀' // U+9C00 <cjk>
	0xEFCE: '鰣' // U+9C23 <cjk>
	0xEFCF: '鱁' // U+9C41 <cjk>
	0xEFD0: '鱏' // U+9C4F <cjk>
	0xEFD1: '鱐' // U+9C50 <cjk>
	0xEFD2: '鱓' // U+9C53 <cjk>
	0xEFD3: '鱣' // U+9C63 <cjk>
	0xEFD4: '鱥' // U+9C65 <cjk>
	0xEFD5: '鱷' // U+9C77 <cjk>
	0xEFD6: '鴝' // U+9D1D <cjk>
	0xEFD7: '鴞' // U+9D1E <cjk>
	0xEFD8: '鵃' // U+9D43 <cjk>
	0xEFD9: '鵇' // U+9D47 <cjk>
	0xEFDA: '鵒' // U+9D52 <cjk>
	0xEFDB: '鵣' // U+9D63 <cjk>
	0xEFDC: '鵰' // U+9D70 <cjk>
	0xEFDD: '鵼' // U+9D7C <cjk>
	0xEFDE: '鶊' // U+9D8A <cjk>
	0xEFDF: '鶖' // U+9D96 <cjk>
	0xEFE0: '鷀' // U+9DC0 <cjk>
	0xEFE1: '鶬' // U+9DAC <cjk>
	0xEFE2: '鶼' // U+9DBC <cjk>
	0xEFE3: '鷗' // U+9DD7 <cjk>
	0xEFE4: '𪆐' // U+2A190 <cjk>
	0xEFE5: '鷧' // U+9DE7 <cjk>
	0xEFE6: '鸇' // U+9E07 <cjk>
	0xEFE7: '鸕' // U+9E15 <cjk>
	0xEFE8: '鹼' // U+9E7C <cjk>
	0xEFE9: '麞' // U+9E9E <cjk>
	0xEFEA: '麤' // U+9EA4 <cjk>
	0xEFEB: '麬' // U+9EAC <cjk>
	0xEFEC: '麯' // U+9EAF <cjk>
	0xEFED: '麴' // U+9EB4 <cjk>
	0xEFEE: '麵' // U+9EB5 <cjk>
	0xEFEF: '黃' // U+9EC3 <cjk>
	0xEFF0: '黑' // U+9ED1 <cjk>
	0xEFF1: '鼐' // U+9F10 <cjk>
	0xEFF2: '鼹' // U+9F39 <cjk>
	0xEFF3: '齗' // U+9F57 <cjk>
	0xEFF4: '龐' // U+9F90 <cjk>
	0xEFF5: '龔' // U+9F94 <cjk>
	0xEFF6: '龗' // U+9F97 <cjk>
	0xEFF7: '龢' // U+9FA2 <cjk>
	0xEFF8: '姸' // U+59F8 <cjk>
	0xEFF9: '屛' // U+5C5B <cjk>
	0xEFFA: '幷' // U+5E77 <cjk>
	0xEFFB: '瘦' // U+7626 <cjk>
	0xEFFC: '繫' // U+7E6B <cjk>
	0xF040: '𠂉' // U+20089 <cjk>
	0xF041: '丂' // U+4E02 <cjk>
	0xF042: '丏' // U+4E0F <cjk>
	0xF043: '丒' // U+4E12 <cjk>
	0xF044: '丩' // U+4E29 <cjk>
	0xF045: '丫' // U+4E2B <cjk>
	0xF046: '丮' // U+4E2E <cjk>
	0xF047: '乀' // U+4E40 <cjk>
	0xF048: '乇' // U+4E47 <cjk>
	0xF049: '么' // U+4E48 <cjk>
	0xF04A: '𠂢' // U+200A2 <cjk>
	0xF04B: '乑' // U+4E51 <cjk>
	0xF04C: '㐆' // U+3406 <cjk>
	0xF04D: '𠂤' // U+200A4 <cjk>
	0xF04E: '乚' // U+4E5A <cjk>
	0xF04F: '乩' // U+4E69 <cjk>
	0xF050: '亝' // U+4E9D <cjk>
	0xF051: '㐬' // U+342C <cjk>
	0xF052: '㐮' // U+342E <cjk>
	0xF053: '亹' // U+4EB9 <cjk>
	0xF054: '亻' // U+4EBB <cjk>
	0xF055: '𠆢' // U+201A2 <cjk>
	0xF056: '亼' // U+4EBC <cjk>
	0xF057: '仃' // U+4EC3 <cjk>
	0xF058: '仈' // U+4EC8 <cjk>
	0xF059: '仐' // U+4ED0 <cjk>
	0xF05A: '仫' // U+4EEB <cjk>
	0xF05B: '仚' // U+4EDA <cjk>
	0xF05C: '仱' // U+4EF1 <cjk>
	0xF05D: '仵' // U+4EF5 <cjk>
	0xF05E: '伀' // U+4F00 <cjk>
	0xF05F: '伖' // U+4F16 <cjk>
	0xF060: '佤' // U+4F64 <cjk>
	0xF061: '伷' // U+4F37 <cjk>
	0xF062: '伾' // U+4F3E <cjk>
	0xF063: '佔' // U+4F54 <cjk>
	0xF064: '佘' // U+4F58 <cjk>
	0xF065: '𠈓' // U+20213 <cjk>
	0xF066: '佷' // U+4F77 <cjk>
	0xF067: '佸' // U+4F78 <cjk>
	0xF068: '佺' // U+4F7A <cjk>
	0xF069: '佽' // U+4F7D <cjk>
	0xF06A: '侂' // U+4F82 <cjk>
	0xF06B: '侅' // U+4F85 <cjk>
	0xF06C: '侒' // U+4F92 <cjk>
	0xF06D: '侚' // U+4F9A <cjk>
	0xF06E: '俦' // U+4FE6 <cjk>
	0xF06F: '侲' // U+4FB2 <cjk>
	0xF070: '侾' // U+4FBE <cjk>
	0xF071: '俅' // U+4FC5 <cjk>
	0xF072: '俋' // U+4FCB <cjk>
	0xF073: '俏' // U+4FCF <cjk>
	0xF074: '俒' // U+4FD2 <cjk>
	0xF075: '㑪' // U+346A <cjk>
	0xF076: '俲' // U+4FF2 <cjk>
	0xF077: '倀' // U+5000 <cjk>
	0xF078: '倐' // U+5010 <cjk>
	0xF079: '倓' // U+5013 <cjk>
	0xF07A: '倜' // U+501C <cjk>
	0xF07B: '倞' // U+501E <cjk>
	0xF07C: '倢' // U+5022 <cjk>
	0xF07D: '㑨' // U+3468 <cjk>
	0xF07E: '偂' // U+5042 <cjk>
	0xF080: '偆' // U+5046 <cjk>
	0xF081: '偎' // U+504E <cjk>
	0xF082: '偓' // U+5053 <cjk>
	0xF083: '偗' // U+5057 <cjk>
	0xF084: '偣' // U+5063 <cjk>
	0xF085: '偦' // U+5066 <cjk>
	0xF086: '偪' // U+506A <cjk>
	0xF087: '偰' // U+5070 <cjk>
	0xF088: '傣' // U+50A3 <cjk>
	0xF089: '傈' // U+5088 <cjk>
	0xF08A: '傒' // U+5092 <cjk>
	0xF08B: '傓' // U+5093 <cjk>
	0xF08C: '傕' // U+5095 <cjk>
	0xF08D: '傖' // U+5096 <cjk>
	0xF08E: '傜' // U+509C <cjk>
	0xF08F: '傪' // U+50AA <cjk>
	0xF090: '𠌫' // U+2032B <cjk>
	0xF091: '傱' // U+50B1 <cjk>
	0xF092: '傺' // U+50BA <cjk>
	0xF093: '傻' // U+50BB <cjk>
	0xF094: '僄' // U+50C4 <cjk>
	0xF095: '僇' // U+50C7 <cjk>
	0xF096: '僳' // U+50F3 <cjk>
	0xF097: '𠎁' // U+20381 <cjk>
	0xF098: '僎' // U+50CE <cjk>
	0xF099: '𠍱' // U+20371 <cjk>
	0xF09A: '僔' // U+50D4 <cjk>
	0xF09B: '僙' // U+50D9 <cjk>
	0xF09C: '僡' // U+50E1 <cjk>
	0xF09D: '僩' // U+50E9 <cjk>
	0xF09E: '㒒' // U+3492 <cjk>
	0xF09F: '宖' // U+5B96 <cjk>
	0xF0A0: '宬' // U+5BAC <cjk>
	0xF0A1: '㝡' // U+3761 <cjk>
	0xF0A2: '寀' // U+5BC0 <cjk>
	0xF0A3: '㝢' // U+3762 <cjk>
	0xF0A4: '寎' // U+5BCE <cjk>
	0xF0A5: '寖' // U+5BD6 <cjk>
	0xF0A6: '㝬' // U+376C <cjk>
	0xF0A7: '㝫' // U+376B <cjk>
	0xF0A8: '寱' // U+5BF1 <cjk>
	0xF0A9: '寽' // U+5BFD <cjk>
	0xF0AA: '㝵' // U+3775 <cjk>
	0xF0AB: '尃' // U+5C03 <cjk>
	0xF0AC: '尩' // U+5C29 <cjk>
	0xF0AD: '尰' // U+5C30 <cjk>
	0xF0AE: '𡱖' // U+21C56 <cjk>
	0xF0AF: '屟' // U+5C5F <cjk>
	0xF0B0: '屣' // U+5C63 <cjk>
	0xF0B1: '屧' // U+5C67 <cjk>
	0xF0B2: '屨' // U+5C68 <cjk>
	0xF0B3: '屩' // U+5C69 <cjk>
	0xF0B4: '屰' // U+5C70 <cjk>
	0xF0B5: '𡴭' // U+21D2D <cjk>
	0xF0B6: '𡵅' // U+21D45 <cjk>
	0xF0B7: '屼' // U+5C7C <cjk>
	0xF0B8: '𡵸' // U+21D78 <cjk>
	0xF0B9: '𡵢' // U+21D62 <cjk>
	0xF0BA: '岈' // U+5C88 <cjk>
	0xF0BB: '岊' // U+5C8A <cjk>
	0xF0BC: '㟁' // U+37C1 <cjk>
	0xF0BD: '𡶡' // U+21DA1 <cjk>
	0xF0BE: '𡶜' // U+21D9C <cjk>
	0xF0BF: '岠' // U+5CA0 <cjk>
	0xF0C0: '岢' // U+5CA2 <cjk>
	0xF0C1: '岦' // U+5CA6 <cjk>
	0xF0C2: '岧' // U+5CA7 <cjk>
	0xF0C3: '𡶒' // U+21D92 <cjk>
	0xF0C4: '岭' // U+5CAD <cjk>
	0xF0C5: '岵' // U+5CB5 <cjk>
	0xF0C6: '𡶷' // U+21DB7 <cjk>
	0xF0C7: '峉' // U+5CC9 <cjk>
	0xF0C8: '𡷠' // U+21DE0 <cjk>
	0xF0C9: '𡸳' // U+21E33 <cjk>
	0xF0CA: '崆' // U+5D06 <cjk>
	0xF0CB: '崐' // U+5D10 <cjk>
	0xF0CC: '崫' // U+5D2B <cjk>
	0xF0CD: '崝' // U+5D1D <cjk>
	0xF0CE: '崠' // U+5D20 <cjk>
	0xF0CF: '崤' // U+5D24 <cjk>
	0xF0D0: '崦' // U+5D26 <cjk>
	0xF0D1: '崱' // U+5D31 <cjk>
	0xF0D2: '崹' // U+5D39 <cjk>
	0xF0D3: '嵂' // U+5D42 <cjk>
	0xF0D4: '㟨' // U+37E8 <cjk>
	0xF0D5: '嵡' // U+5D61 <cjk>
	0xF0D6: '嵪' // U+5D6A <cjk>
	0xF0D7: '㟴' // U+37F4 <cjk>
	0xF0D8: '嵰' // U+5D70 <cjk>
	0xF0D9: '𡼞' // U+21F1E <cjk>
	0xF0DA: '㟽' // U+37FD <cjk>
	0xF0DB: '嶈' // U+5D88 <cjk>
	0xF0DC: '㠀' // U+3800 <cjk>
	0xF0DD: '嶒' // U+5D92 <cjk>
	0xF0DE: '嶔' // U+5D94 <cjk>
	0xF0DF: '嶗' // U+5D97 <cjk>
	0xF0E0: '嶙' // U+5D99 <cjk>
	0xF0E1: '嶰' // U+5DB0 <cjk>
	0xF0E2: '嶲' // U+5DB2 <cjk>
	0xF0E3: '嶴' // U+5DB4 <cjk>
	0xF0E4: '𡽶' // U+21F76 <cjk>
	0xF0E5: '嶹' // U+5DB9 <cjk>
	0xF0E6: '巑' // U+5DD1 <cjk>
	0xF0E7: '巗' // U+5DD7 <cjk>
	0xF0E8: '巘' // U+5DD8 <cjk>
	0xF0E9: '巠' // U+5DE0 <cjk>
	0xF0EA: '𡿺' // U+21FFA <cjk>
	0xF0EB: '巤' // U+5DE4 <cjk>
	0xF0EC: '巩' // U+5DE9 <cjk>
	0xF0ED: '㠯' // U+382F <cjk>
	0xF0EE: '帀' // U+5E00 <cjk>
	0xF0EF: '㠶' // U+3836 <cjk>
	0xF0F0: '帒' // U+5E12 <cjk>
	0xF0F1: '帕' // U+5E15 <cjk>
	0xF0F2: '㡀' // U+3840 <cjk>
	0xF0F3: '帟' // U+5E1F <cjk>
	0xF0F4: '帮' // U+5E2E <cjk>
	0xF0F5: '帾' // U+5E3E <cjk>
	0xF0F6: '幉' // U+5E49 <cjk>
	0xF0F7: '㡜' // U+385C <cjk>
	0xF0F8: '幖' // U+5E56 <cjk>
	0xF0F9: '㡡' // U+3861 <cjk>
	0xF0FA: '幫' // U+5E6B <cjk>
	0xF0FB: '幬' // U+5E6C <cjk>
	0xF0FC: '幭' // U+5E6D <cjk>
	0xF140: '儈' // U+5108 <cjk>
	0xF141: '𠏹' // U+203F9 <cjk>
	0xF142: '儗' // U+5117 <cjk>
	0xF143: '儛' // U+511B <cjk>
	0xF144: '𠑊' // U+2044A <cjk>
	0xF145: '兠' // U+5160 <cjk>
	0xF146: '𠔉' // U+20509 <cjk>
	0xF147: '关' // U+5173 <cjk>
	0xF148: '冃' // U+5183 <cjk>
	0xF149: '冋' // U+518B <cjk>
	0xF14A: '㒼' // U+34BC <cjk>
	0xF14B: '冘' // U+5198 <cjk>
	0xF14C: '冣' // U+51A3 <cjk>
	0xF14D: '冭' // U+51AD <cjk>
	0xF14E: '㓇' // U+34C7 <cjk>
	0xF14F: '冼' // U+51BC <cjk>
	0xF150: '𠗖' // U+205D6 <cjk>
	0xF151: '𠘨' // U+20628 <cjk>
	0xF152: '凳' // U+51F3 <cjk>
	0xF153: '凴' // U+51F4 <cjk>
	0xF154: '刂' // U+5202 <cjk>
	0xF155: '划' // U+5212 <cjk>
	0xF156: '刖' // U+5216 <cjk>
	0xF157: '𠝏' // U+2074F <cjk>
	0xF158: '剕' // U+5255 <cjk>
	0xF159: '剜' // U+525C <cjk>
	0xF15A: '剬' // U+526C <cjk>
	0xF15B: '剷' // U+5277 <cjk>
	0xF15C: '劄' // U+5284 <cjk>
	0xF15D: '劂' // U+5282 <cjk>
	0xF15E: '𠠇' // U+20807 <cjk>
	0xF15F: '劘' // U+5298 <cjk>
	0xF160: '𠠺' // U+2083A <cjk>
	0xF161: '劤' // U+52A4 <cjk>
	0xF162: '劦' // U+52A6 <cjk>
	0xF163: '劯' // U+52AF <cjk>
	0xF164: '劺' // U+52BA <cjk>
	0xF165: '劻' // U+52BB <cjk>
	0xF166: '勊' // U+52CA <cjk>
	0xF167: '㔟' // U+351F <cjk>
	0xF168: '勑' // U+52D1 <cjk>
	0xF169: '𠢹' // U+208B9 <cjk>
	0xF16A: '勷' // U+52F7 <cjk>
	0xF16B: '匊' // U+530A <cjk>
	0xF16C: '匋' // U+530B <cjk>
	0xF16D: '匤' // U+5324 <cjk>
	0xF16E: '匵' // U+5335 <cjk>
	0xF16F: '匾' // U+533E <cjk>
	0xF170: '卂' // U+5342 <cjk>
	0xF171: '𠥼' // U+2097C <cjk>
	0xF172: '𠦝' // U+2099D <cjk>
	0xF173: '卧' // U+5367 <cjk>
	0xF174: '卬' // U+536C <cjk>
	0xF175: '卺' // U+537A <cjk>
	0xF176: '厤' // U+53A4 <cjk>
	0xF177: '厴' // U+53B4 <cjk>
	0xF178: '𠫓' // U+20AD3 <cjk>
	0xF179: '厷' // U+53B7 <cjk>
	0xF17A: '叀' // U+53C0 <cjk>
	0xF17B: '𠬝' // U+20B1D <cjk>
	0xF17C: '㕝' // U+355D <cjk>
	0xF17D: '㕞' // U+355E <cjk>
	0xF17E: '叕' // U+53D5 <cjk>
	0xF180: '叚' // U+53DA <cjk>
	0xF181: '㕣' // U+3563 <cjk>
	0xF182: '叴' // U+53F4 <cjk>
	0xF183: '叵' // U+53F5 <cjk>
	0xF184: '呕' // U+5455 <cjk>
	0xF185: '吤' // U+5424 <cjk>
	0xF186: '吨' // U+5428 <cjk>
	0xF187: '㕮' // U+356E <cjk>
	0xF188: '呃' // U+5443 <cjk>
	0xF189: '呢' // U+5462 <cjk>
	0xF18A: '呦' // U+5466 <cjk>
	0xF18B: '呬' // U+546C <cjk>
	0xF18C: '咊' // U+548A <cjk>
	0xF18D: '咍' // U+548D <cjk>
	0xF18E: '咕' // U+5495 <cjk>
	0xF18F: '咠' // U+54A0 <cjk>
	0xF190: '咦' // U+54A6 <cjk>
	0xF191: '咭' // U+54AD <cjk>
	0xF192: '咮' // U+54AE <cjk>
	0xF193: '咷' // U+54B7 <cjk>
	0xF194: '咺' // U+54BA <cjk>
	0xF195: '咿' // U+54BF <cjk>
	0xF196: '哃' // U+54C3 <cjk>
	0xF197: '𠵅' // U+20D45 <cjk>
	0xF198: '哬' // U+54EC <cjk>
	0xF199: '哯' // U+54EF <cjk>
	0xF19A: '哱' // U+54F1 <cjk>
	0xF19B: '哳' // U+54F3 <cjk>
	0xF19C: '唀' // U+5500 <cjk>
	0xF19D: '唁' // U+5501 <cjk>
	0xF19E: '唉' // U+5509 <cjk>
	0xF19F: '唼' // U+553C <cjk>
	0xF1A0: '啁' // U+5541 <cjk>
	0xF1A1: '㖦' // U+35A6 <cjk>
	0xF1A2: '啇' // U+5547 <cjk>
	0xF1A3: '啊' // U+554A <cjk>
	0xF1A4: '㖨' // U+35A8 <cjk>
	0xF1A5: '啠' // U+5560 <cjk>
	0xF1A6: '啡' // U+5561 <cjk>
	0xF1A7: '啤' // U+5564 <cjk>
	0xF1A8: '𠷡' // U+20DE1 <cjk>
	0xF1A9: '啽' // U+557D <cjk>
	0xF1AA: '喂' // U+5582 <cjk>
	0xF1AB: '喈' // U+5588 <cjk>
	0xF1AC: '喑' // U+5591 <cjk>
	0xF1AD: '㗅' // U+35C5 <cjk>
	0xF1AE: '嗒' // U+55D2 <cjk>
	0xF1AF: '𠺕' // U+20E95 <cjk>
	0xF1B0: '𠹭' // U+20E6D <cjk>
	0xF1B1: '喿' // U+55BF <cjk>
	0xF1B2: '嗉' // U+55C9 <cjk>
	0xF1B3: '嗌' // U+55CC <cjk>
	0xF1B4: '嗑' // U+55D1 <cjk>
	0xF1B5: '嗝' // U+55DD <cjk>
	0xF1B6: '㗚' // U+35DA <cjk>
	0xF1B7: '嗢' // U+55E2 <cjk>
	0xF1B8: '𠹤' // U+20E64 <cjk>
	0xF1B9: '嗩' // U+55E9 <cjk>
	0xF1BA: '嘨' // U+5628 <cjk>
	0xF1BB: '𠽟' // U+20F5F <cjk>
	0xF1BC: '嘇' // U+5607 <cjk>
	0xF1BD: '嘐' // U+5610 <cjk>
	0xF1BE: '嘰' // U+5630 <cjk>
	0xF1BF: '嘷' // U+5637 <cjk>
	0xF1C0: '㗴' // U+35F4 <cjk>
	0xF1C1: '嘽' // U+563D <cjk>
	0xF1C2: '嘿' // U+563F <cjk>
	0xF1C3: '噀' // U+5640 <cjk>
	0xF1C4: '噇' // U+5647 <cjk>
	0xF1C5: '噞' // U+565E <cjk>
	0xF1C6: '噠' // U+5660 <cjk>
	0xF1C7: '噭' // U+566D <cjk>
	0xF1C8: '㘅' // U+3605 <cjk>
	0xF1C9: '嚈' // U+5688 <cjk>
	0xF1CA: '嚌' // U+568C <cjk>
	0xF1CB: '嚕' // U+5695 <cjk>
	0xF1CC: '嚚' // U+569A <cjk>
	0xF1CD: '嚝' // U+569D <cjk>
	0xF1CE: '嚨' // U+56A8 <cjk>
	0xF1CF: '嚭' // U+56AD <cjk>
	0xF1D0: '嚲' // U+56B2 <cjk>
	0xF1D1: '囅' // U+56C5 <cjk>
	0xF1D2: '囍' // U+56CD <cjk>
	0xF1D3: '囟' // U+56DF <cjk>
	0xF1D4: '囨' // U+56E8 <cjk>
	0xF1D5: '囶' // U+56F6 <cjk>
	0xF1D6: '囷' // U+56F7 <cjk>
	0xF1D7: '𡈁' // U+21201 <cjk>
	0xF1D8: '圕' // U+5715 <cjk>
	0xF1D9: '圣' // U+5723 <cjk>
	0xF1DA: '𡉕' // U+21255 <cjk>
	0xF1DB: '圩' // U+5729 <cjk>
	0xF1DC: '𡉻' // U+2127B <cjk>
	0xF1DD: '坅' // U+5745 <cjk>
	0xF1DE: '坆' // U+5746 <cjk>
	0xF1DF: '坌' // U+574C <cjk>
	0xF1E0: '坍' // U+574D <cjk>
	0xF1E1: '𡉴' // U+21274 <cjk>
	0xF1E2: '坨' // U+5768 <cjk>
	0xF1E3: '坯' // U+576F <cjk>
	0xF1E4: '坳' // U+5773 <cjk>
	0xF1E5: '坴' // U+5774 <cjk>
	0xF1E6: '坵' // U+5775 <cjk>
	0xF1E7: '坻' // U+577B <cjk>
	0xF1E8: '𡋤' // U+212E4 <cjk>
	0xF1E9: '𡋗' // U+212D7 <cjk>
	0xF1EA: '垬' // U+57AC <cjk>
	0xF1EB: '垚' // U+579A <cjk>
	0xF1EC: '垝' // U+579D <cjk>
	0xF1ED: '垞' // U+579E <cjk>
	0xF1EE: '垨' // U+57A8 <cjk>
	0xF1EF: '埗' // U+57D7 <cjk>
	0xF1F0: '𡋽' // U+212FD <cjk>
	0xF1F1: '埌' // U+57CC <cjk>
	0xF1F2: '𡌶' // U+21336 <cjk>
	0xF1F3: '𡍄' // U+21344 <cjk>
	0xF1F4: '埞' // U+57DE <cjk>
	0xF1F5: '埦' // U+57E6 <cjk>
	0xF1F6: '埰' // U+57F0 <cjk>
	0xF1F7: '㙊' // U+364A <cjk>
	0xF1F8: '埸' // U+57F8 <cjk>
	0xF1F9: '埻' // U+57FB <cjk>
	0xF1FA: '埽' // U+57FD <cjk>
	0xF1FB: '堄' // U+5804 <cjk>
	0xF1FC: '堞' // U+581E <cjk>
	0xF240: '堠' // U+5820 <cjk>
	0xF241: '堧' // U+5827 <cjk>
	0xF242: '堲' // U+5832 <cjk>
	0xF243: '堹' // U+5839 <cjk>
	0xF244: '𡏄' // U+213C4 <cjk>
	0xF245: '塉' // U+5849 <cjk>
	0xF246: '塌' // U+584C <cjk>
	0xF247: '塧' // U+5867 <cjk>
	0xF248: '墊' // U+588A <cjk>
	0xF249: '墋' // U+588B <cjk>
	0xF24A: '墍' // U+588D <cjk>
	0xF24B: '墏' // U+588F <cjk>
	0xF24C: '墐' // U+5890 <cjk>
	0xF24D: '墔' // U+5894 <cjk>
	0xF24E: '墝' // U+589D <cjk>
	0xF24F: '墪' // U+58AA <cjk>
	0xF250: '墱' // U+58B1 <cjk>
	0xF251: '𡑭' // U+2146D <cjk>
	0xF252: '壃' // U+58C3 <cjk>
	0xF253: '壍' // U+58CD <cjk>
	0xF254: '壢' // U+58E2 <cjk>
	0xF255: '壳' // U+58F3 <cjk>
	0xF256: '壴' // U+58F4 <cjk>
	0xF257: '夅' // U+5905 <cjk>
	0xF258: '夆' // U+5906 <cjk>
	0xF259: '夋' // U+590B <cjk>
	0xF25A: '复' // U+590D <cjk>
	0xF25B: '夔' // U+5914 <cjk>
	0xF25C: '夤' // U+5924 <cjk>
	0xF25D: '𡗗' // U+215D7 <cjk>
	0xF25E: '㚑' // U+3691 <cjk>
	0xF25F: '夽' // U+593D <cjk>
	0xF260: '㚙' // U+3699 <cjk>
	0xF261: '奆' // U+5946 <cjk>
	0xF262: '㚖' // U+3696 <cjk>
	0xF263: '𦰩' // U+26C29 <cjk>
	0xF264: '奛' // U+595B <cjk>
	0xF265: '奟' // U+595F <cjk>
	0xF266: '𡙇' // U+21647 <cjk>
	0xF267: '奵' // U+5975 <cjk>
	0xF268: '奶' // U+5976 <cjk>
	0xF269: '奼' // U+597C <cjk>
	0xF26A: '妟' // U+599F <cjk>
	0xF26B: '妮' // U+59AE <cjk>
	0xF26C: '妼' // U+59BC <cjk>
	0xF26D: '姈' // U+59C8 <cjk>
	0xF26E: '姍' // U+59CD <cjk>
	0xF26F: '姞' // U+59DE <cjk>
	0xF270: '姣' // U+59E3 <cjk>
	0xF271: '姤' // U+59E4 <cjk>
	0xF272: '姧' // U+59E7 <cjk>
	0xF273: '姮' // U+59EE <cjk>
	0xF274: '𡜆' // U+21706 <cjk>
	0xF275: '𡝂' // U+21742 <cjk>
	0xF276: '㛏' // U+36CF <cjk>
	0xF277: '娌' // U+5A0C <cjk>
	0xF278: '娍' // U+5A0D <cjk>
	0xF279: '娗' // U+5A17 <cjk>
	0xF27A: '娧' // U+5A27 <cjk>
	0xF27B: '娭' // U+5A2D <cjk>
	0xF27C: '婕' // U+5A55 <cjk>
	0xF27D: '婥' // U+5A65 <cjk>
	0xF27E: '婺' // U+5A7A <cjk>
	0xF280: '媋' // U+5A8B <cjk>
	0xF281: '媜' // U+5A9C <cjk>
	0xF282: '媟' // U+5A9F <cjk>
	0xF283: '媠' // U+5AA0 <cjk>
	0xF284: '媢' // U+5AA2 <cjk>
	0xF285: '媱' // U+5AB1 <cjk>
	0xF286: '媳' // U+5AB3 <cjk>
	0xF287: '媵' // U+5AB5 <cjk>
	0xF288: '媺' // U+5ABA <cjk>
	0xF289: '媿' // U+5ABF <cjk>
	0xF28A: '嫚' // U+5ADA <cjk>
	0xF28B: '嫜' // U+5ADC <cjk>
	0xF28C: '嫠' // U+5AE0 <cjk>
	0xF28D: '嫥' // U+5AE5 <cjk>
	0xF28E: '嫰' // U+5AF0 <cjk>
	0xF28F: '嫮' // U+5AEE <cjk>
	0xF290: '嫵' // U+5AF5 <cjk>
	0xF291: '嬀' // U+5B00 <cjk>
	0xF292: '嬈' // U+5B08 <cjk>
	0xF293: '嬗' // U+5B17 <cjk>
	0xF294: '嬴' // U+5B34 <cjk>
	0xF295: '嬭' // U+5B2D <cjk>
	0xF296: '孌' // U+5B4C <cjk>
	0xF297: '孒' // U+5B52 <cjk>
	0xF298: '孨' // U+5B68 <cjk>
	0xF299: '孯' // U+5B6F <cjk>
	0xF29A: '孼' // U+5B7C <cjk>
	0xF29B: '孿' // U+5B7F <cjk>
	0xF29C: '宁' // U+5B81 <cjk>
	0xF29D: '宄' // U+5B84 <cjk>
	0xF29E: '𡧃' // U+219C3 <cjk>
	0xF29F: '幮' // U+5E6E <cjk>
	0xF2A0: '𢅻' // U+2217B <cjk>
	0xF2A1: '庥' // U+5EA5 <cjk>
	0xF2A2: '庪' // U+5EAA <cjk>
	0xF2A3: '庬' // U+5EAC <cjk>
	0xF2A4: '庹' // U+5EB9 <cjk>
	0xF2A5: '庿' // U+5EBF <cjk>
	0xF2A6: '廆' // U+5EC6 <cjk>
	0xF2A7: '廒' // U+5ED2 <cjk>
	0xF2A8: '廙' // U+5ED9 <cjk>
	0xF2A9: '𢌞' // U+2231E <cjk>
	0xF2AA: '廽' // U+5EFD <cjk>
	0xF2AB: '弈' // U+5F08 <cjk>
	0xF2AC: '弎' // U+5F0E <cjk>
	0xF2AD: '弜' // U+5F1C <cjk>
	0xF2AE: '𢎭' // U+223AD <cjk>
	0xF2AF: '弞' // U+5F1E <cjk>
	0xF2B0: '彇' // U+5F47 <cjk>
	0xF2B1: '彣' // U+5F63 <cjk>
	0xF2B2: '彲' // U+5F72 <cjk>
	0xF2B3: '彾' // U+5F7E <cjk>
	0xF2B4: '徏' // U+5F8F <cjk>
	0xF2B5: '徢' // U+5FA2 <cjk>
	0xF2B6: '徤' // U+5FA4 <cjk>
	0xF2B7: '徸' // U+5FB8 <cjk>
	0xF2B8: '忄' // U+5FC4 <cjk>
	0xF2B9: '㣺' // U+38FA <cjk>
	0xF2BA: '忇' // U+5FC7 <cjk>
	0xF2BB: '忋' // U+5FCB <cjk>
	0xF2BC: '忒' // U+5FD2 <cjk>
	0xF2BD: '忓' // U+5FD3 <cjk>
	0xF2BE: '忔' // U+5FD4 <cjk>
	0xF2BF: '忢' // U+5FE2 <cjk>
	0xF2C0: '忮' // U+5FEE <cjk>
	0xF2C1: '忯' // U+5FEF <cjk>
	0xF2C2: '忳' // U+5FF3 <cjk>
	0xF2C3: '忼' // U+5FFC <cjk>
	0xF2C4: '㤗' // U+3917 <cjk>
	0xF2C5: '怗' // U+6017 <cjk>
	0xF2C6: '怢' // U+6022 <cjk>
	0xF2C7: '怤' // U+6024 <cjk>
	0xF2C8: '㤚' // U+391A <cjk>
	0xF2C9: '恌' // U+604C <cjk>
	0xF2CA: '恿' // U+607F <cjk>
	0xF2CB: '悊' // U+608A <cjk>
	0xF2CC: '悕' // U+6095 <cjk>
	0xF2CD: '您' // U+60A8 <cjk>
	0xF2CE: '𢛳' // U+226F3 <cjk>
	0xF2CF: '悰' // U+60B0 <cjk>
	0xF2D0: '悱' // U+60B1 <cjk>
	0xF2D1: '悾' // U+60BE <cjk>
	0xF2D2: '惈' // U+60C8 <cjk>
	0xF2D3: '惙' // U+60D9 <cjk>
	0xF2D4: '惛' // U+60DB <cjk>
	0xF2D5: '惮' // U+60EE <cjk>
	0xF2D6: '惲' // U+60F2 <cjk>
	0xF2D7: '惵' // U+60F5 <cjk>
	0xF2D8: '愐' // U+6110 <cjk>
	0xF2D9: '愒' // U+6112 <cjk>
	0xF2DA: '愓' // U+6113 <cjk>
	0xF2DB: '愙' // U+6119 <cjk>
	0xF2DC: '愞' // U+611E <cjk>
	0xF2DD: '愺' // U+613A <cjk>
	0xF2DE: '㥯' // U+396F <cjk>
	0xF2DF: '慁' // U+6141 <cjk>
	0xF2E0: '慆' // U+6146 <cjk>
	0xF2E1: '慠' // U+6160 <cjk>
	0xF2E2: '慼' // U+617C <cjk>
	0xF2E3: '𢡛' // U+2285B <cjk>
	0xF2E4: '憒' // U+6192 <cjk>
	0xF2E5: '憓' // U+6193 <cjk>
	0xF2E6: '憗' // U+6197 <cjk>
	0xF2E7: '憘' // U+6198 <cjk>
	0xF2E8: '憥' // U+61A5 <cjk>
	0xF2E9: '憨' // U+61A8 <cjk>
	0xF2EA: '憭' // U+61AD <cjk>
	0xF2EB: '𢢫' // U+228AB <cjk>
	0xF2EC: '懕' // U+61D5 <cjk>
	0xF2ED: '懝' // U+61DD <cjk>
	0xF2EE: '懟' // U+61DF <cjk>
	0xF2EF: '懵' // U+61F5 <cjk>
	0xF2F0: '𢦏' // U+2298F <cjk>
	0xF2F1: '戕' // U+6215 <cjk>
	0xF2F2: '戣' // U+6223 <cjk>
	0xF2F3: '戩' // U+6229 <cjk>
	0xF2F4: '扆' // U+6246 <cjk>
	0xF2F5: '扌' // U+624C <cjk>
	0xF2F6: '扑' // U+6251 <cjk>
	0xF2F7: '扒' // U+6252 <cjk>
	0xF2F8: '扡' // U+6261 <cjk>
	0xF2F9: '扤' // U+6264 <cjk>
	0xF2FA: '扻' // U+627B <cjk>
	0xF2FB: '扭' // U+626D <cjk>
	0xF2FC: '扳' // U+6273 <cjk>
	0xF340: '抙' // U+6299 <cjk>
	0xF341: '抦' // U+62A6 <cjk>
	0xF342: '拕' // U+62D5 <cjk>
	0xF343: '𢪸' // U+22AB8 <cjk>
	0xF344: '拽' // U+62FD <cjk>
	0xF345: '挃' // U+6303 <cjk>
	0xF346: '挍' // U+630D <cjk>
	0xF347: '挐' // U+6310 <cjk>
	0xF348: '𢭏' // U+22B4F <cjk>
	0xF349: '𢭐' // U+22B50 <cjk>
	0xF34A: '挲' // U+6332 <cjk>
	0xF34B: '挵' // U+6335 <cjk>
	0xF34C: '挻' // U+633B <cjk>
	0xF34D: '挼' // U+633C <cjk>
	0xF34E: '捁' // U+6341 <cjk>
	0xF34F: '捄' // U+6344 <cjk>
	0xF350: '捎' // U+634E <cjk>
	0xF351: '𢭆' // U+22B46 <cjk>
	0xF352: '捙' // U+6359 <cjk>
	0xF353: '𢰝' // U+22C1D <cjk>
	0xF354: '𢮦' // U+22BA6 <cjk>
	0xF355: '捬' // U+636C <cjk>
	0xF356: '掄' // U+6384 <cjk>
	0xF357: '掙' // U+6399 <cjk>
	0xF358: '𢰤' // U+22C24 <cjk>
	0xF359: '掔' // U+6394 <cjk>
	0xF35A: '掽' // U+63BD <cjk>
	0xF35B: '揷' // U+63F7 <cjk>
	0xF35C: '揔' // U+63D4 <cjk>
	0xF35D: '揕' // U+63D5 <cjk>
	0xF35E: '揜' // U+63DC <cjk>
	0xF35F: '揠' // U+63E0 <cjk>
	0xF360: '揫' // U+63EB <cjk>
	0xF361: '揬' // U+63EC <cjk>
	0xF362: '揲' // U+63F2 <cjk>
	0xF363: '搉' // U+6409 <cjk>
	0xF364: '搞' // U+641E <cjk>
	0xF365: '搥' // U+6425 <cjk>
	0xF366: '搩' // U+6429 <cjk>
	0xF367: '搯' // U+642F <cjk>
	0xF368: '摚' // U+645A <cjk>
	0xF369: '摛' // U+645B <cjk>
	0xF36A: '摝' // U+645D <cjk>
	0xF36B: '摳' // U+6473 <cjk>
	0xF36C: '摽' // U+647D <cjk>
	0xF36D: '撇' // U+6487 <cjk>
	0xF36E: '撑' // U+6491 <cjk>
	0xF36F: '撝' // U+649D <cjk>
	0xF370: '撟' // U+649F <cjk>
	0xF371: '擋' // U+64CB <cjk>
	0xF372: '擌' // U+64CC <cjk>
	0xF373: '擕' // U+64D5 <cjk>
	0xF374: '擗' // U+64D7 <cjk>
	0xF375: '𢷡' // U+22DE1 <cjk>
	0xF376: '擤' // U+64E4 <cjk>
	0xF377: '擥' // U+64E5 <cjk>
	0xF378: '擿' // U+64FF <cjk>
	0xF379: '攄' // U+6504 <cjk>
	0xF37A: '㩮' // U+3A6E <cjk>
	0xF37B: '攏' // U+650F <cjk>
	0xF37C: '攔' // U+6514 <cjk>
	0xF37D: '攖' // U+6516 <cjk>
	0xF37E: '㩳' // U+3A73 <cjk>
	0xF380: '攞' // U+651E <cjk>
	0xF381: '攲' // U+6532 <cjk>
	0xF382: '敄' // U+6544 <cjk>
	0xF383: '敔' // U+6554 <cjk>
	0xF384: '敫' // U+656B <cjk>
	0xF385: '敺' // U+657A <cjk>
	0xF386: '斁' // U+6581 <cjk>
	0xF387: '斄' // U+6584 <cjk>
	0xF388: '斅' // U+6585 <cjk>
	0xF389: '斊' // U+658A <cjk>
	0xF38A: '斲' // U+65B2 <cjk>
	0xF38B: '斵' // U+65B5 <cjk>
	0xF38C: '斸' // U+65B8 <cjk>
	0xF38D: '斿' // U+65BF <cjk>
	0xF38E: '旂' // U+65C2 <cjk>
	0xF38F: '旉' // U+65C9 <cjk>
	0xF390: '旔' // U+65D4 <cjk>
	0xF391: '㫖' // U+3AD6 <cjk>
	0xF392: '旲' // U+65F2 <cjk>
	0xF393: '旹' // U+65F9 <cjk>
	0xF394: '旼' // U+65FC <cjk>
	0xF395: '昄' // U+6604 <cjk>
	0xF396: '昈' // U+6608 <cjk>
	0xF397: '昡' // U+6621 <cjk>
	0xF398: '昪' // U+662A <cjk>
	0xF399: '晅' // U+6645 <cjk>
	0xF39A: '晑' // U+6651 <cjk>
	0xF39B: '晎' // U+664E <cjk>
	0xF39C: '㫪' // U+3AEA <cjk>
	0xF39D: '𣇃' // U+231C3 <cjk>
	0xF39E: '晗' // U+6657 <cjk>
	0xF39F: '晛' // U+665B <cjk>
	0xF3A0: '晣' // U+6663 <cjk>
	0xF3A1: '𣇵' // U+231F5 <cjk>
	0xF3A2: '𣆶' // U+231B6 <cjk>
	0xF3A3: '晪' // U+666A <cjk>
	0xF3A4: '晫' // U+666B <cjk>
	0xF3A5: '晬' // U+666C <cjk>
	0xF3A6: '晭' // U+666D <cjk>
	0xF3A7: '晻' // U+667B <cjk>
	0xF3A8: '暀' // U+6680 <cjk>
	0xF3A9: '暐' // U+6690 <cjk>
	0xF3AA: '暒' // U+6692 <cjk>
	0xF3AB: '暙' // U+6699 <cjk>
	0xF3AC: '㬎' // U+3B0E <cjk>
	0xF3AD: '暭' // U+66AD <cjk>
	0xF3AE: '暱' // U+66B1 <cjk>
	0xF3AF: '暵' // U+66B5 <cjk>
	0xF3B0: '㬚' // U+3B1A <cjk>
	0xF3B1: '暿' // U+66BF <cjk>
	0xF3B2: '㬜' // U+3B1C <cjk>
	0xF3B3: '曬' // U+66EC <cjk>
	0xF3B4: '㫗' // U+3AD7 <cjk>
	0xF3B5: '朁' // U+6701 <cjk>
	0xF3B6: '朅' // U+6705 <cjk>
	0xF3B7: '朒' // U+6712 <cjk>
	0xF3B8: '𣍲' // U+23372 <cjk>
	0xF3B9: '朙' // U+6719 <cjk>
	0xF3BA: '𣏓' // U+233D3 <cjk>
	0xF3BB: '𣏒' // U+233D2 <cjk>
	0xF3BC: '杌' // U+674C <cjk>
	0xF3BD: '杍' // U+674D <cjk>
	0xF3BE: '杔' // U+6754 <cjk>
	0xF3BF: '杝' // U+675D <cjk>
	0xF3C0: '𣏐' // U+233D0 <cjk>
	0xF3C1: '𣏤' // U+233E4 <cjk>
	0xF3C2: '𣏕' // U+233D5 <cjk>
	0xF3C3: '杴' // U+6774 <cjk>
	0xF3C4: '杶' // U+6776 <cjk>
	0xF3C5: '𣏚' // U+233DA <cjk>
	0xF3C6: '枒' // U+6792 <cjk>
	0xF3C7: '𣏟' // U+233DF <cjk>
	0xF3C8: '荣' // U+8363 <cjk>
	0xF3C9: '栐' // U+6810 <cjk>
	0xF3CA: '枰' // U+67B0 <cjk>
	0xF3CB: '枲' // U+67B2 <cjk>
	0xF3CC: '柃' // U+67C3 <cjk>
	0xF3CD: '柈' // U+67C8 <cjk>
	0xF3CE: '柒' // U+67D2 <cjk>
	0xF3CF: '柙' // U+67D9 <cjk>
	0xF3D0: '柛' // U+67DB <cjk>
	0xF3D1: '柰' // U+67F0 <cjk>
	0xF3D2: '柷' // U+67F7 <cjk>
	0xF3D3: '𣑊' // U+2344A <cjk>
	0xF3D4: '𣑑' // U+23451 <cjk>
	0xF3D5: '𣑋' // U+2344B <cjk>
	0xF3D6: '栘' // U+6818 <cjk>
	0xF3D7: '栟' // U+681F <cjk>
	0xF3D8: '栭' // U+682D <cjk>
	0xF3D9: '𣑥' // U+23465 <cjk>
	0xF3DA: '栳' // U+6833 <cjk>
	0xF3DB: '栻' // U+683B <cjk>
	0xF3DC: '栾' // U+683E <cjk>
	0xF3DD: '桄' // U+6844 <cjk>
	0xF3DE: '桅' // U+6845 <cjk>
	0xF3DF: '桉' // U+6849 <cjk>
	0xF3E0: '桌' // U+684C <cjk>
	0xF3E1: '桕' // U+6855 <cjk>
	0xF3E2: '桗' // U+6857 <cjk>
	0xF3E3: '㭷' // U+3B77 <cjk>
	0xF3E4: '桫' // U+686B <cjk>
	0xF3E5: '桮' // U+686E <cjk>
	0xF3E6: '桺' // U+687A <cjk>
	0xF3E7: '桼' // U+687C <cjk>
	0xF3E8: '梂' // U+6882 <cjk>
	0xF3E9: '梐' // U+6890 <cjk>
	0xF3EA: '梖' // U+6896 <cjk>
	0xF3EB: '㭭' // U+3B6D <cjk>
	0xF3EC: '梘' // U+6898 <cjk>
	0xF3ED: '梙' // U+6899 <cjk>
	0xF3EE: '梚' // U+689A <cjk>
	0xF3EF: '梜' // U+689C <cjk>
	0xF3F0: '梪' // U+68AA <cjk>
	0xF3F1: '梫' // U+68AB <cjk>
	0xF3F2: '梴' // U+68B4 <cjk>
	0xF3F3: '梻' // U+68BB <cjk>
	0xF3F4: '棻' // U+68FB <cjk>
	0xF3F5: '𣓤' // U+234E4 <cjk>
	0xF3F6: '𣕚' // U+2355A <cjk>
	0xF3F7: '﨓' // U+FA13 CJK COMPATIBILITY IDEOGRAPH-FA13
	0xF3F8: '棃' // U+68C3 <cjk>
	0xF3F9: '棅' // U+68C5 <cjk>
	0xF3FA: '棌' // U+68CC <cjk>
	0xF3FB: '棏' // U+68CF <cjk>
	0xF3FC: '棖' // U+68D6 <cjk>
	0xF440: '棙' // U+68D9 <cjk>
	0xF441: '棤' // U+68E4 <cjk>
	0xF442: '棥' // U+68E5 <cjk>
	0xF443: '棬' // U+68EC <cjk>
	0xF444: '棷' // U+68F7 <cjk>
	0xF445: '椃' // U+6903 <cjk>
	0xF446: '椇' // U+6907 <cjk>
	0xF447: '㮇' // U+3B87 <cjk>
	0xF448: '㮈' // U+3B88 <cjk>
	0xF449: '𣖔' // U+23594 <cjk>
	0xF44A: '椻' // U+693B <cjk>
	0xF44B: '㮍' // U+3B8D <cjk>
	0xF44C: '楆' // U+6946 <cjk>
	0xF44D: '楩' // U+6969 <cjk>
	0xF44E: '楬' // U+696C <cjk>
	0xF44F: '楲' // U+6972 <cjk>
	0xF450: '楺' // U+697A <cjk>
	0xF451: '楿' // U+697F <cjk>
	0xF452: '榒' // U+6992 <cjk>
	0xF453: '㮤' // U+3BA4 <cjk>
	0xF454: '榖' // U+6996 <cjk>
	0xF455: '榘' // U+6998 <cjk>
	0xF456: '榦' // U+69A6 <cjk>
	0xF457: '榰' // U+69B0 <cjk>
	0xF458: '榷' // U+69B7 <cjk>
	0xF459: '榺' // U+69BA <cjk>
	0xF45A: '榼' // U+69BC <cjk>
	0xF45B: '槀' // U+69C0 <cjk>
	0xF45C: '槑' // U+69D1 <cjk>
	0xF45D: '槖' // U+69D6 <cjk>
	0xF45E: '𣘹' // U+23639 <cjk>
	0xF45F: '𣙇' // U+23647 <cjk>
	0xF460: '樰' // U+6A30 <cjk>
	0xF461: '𣘸' // U+23638 <cjk>
	0xF462: '𣘺' // U+2363A <cjk>
	0xF463: '槣' // U+69E3 <cjk>
	0xF464: '槮' // U+69EE <cjk>
	0xF465: '槯' // U+69EF <cjk>
	0xF466: '槳' // U+69F3 <cjk>
	0xF467: '㯍' // U+3BCD <cjk>
	0xF468: '槴' // U+69F4 <cjk>
	0xF469: '槾' // U+69FE <cjk>
	0xF46A: '樑' // U+6A11 <cjk>
	0xF46B: '樚' // U+6A1A <cjk>
	0xF46C: '樝' // U+6A1D <cjk>
	0xF46D: '𣜜' // U+2371C <cjk>
	0xF46E: '樲' // U+6A32 <cjk>
	0xF46F: '樳' // U+6A33 <cjk>
	0xF470: '樴' // U+6A34 <cjk>
	0xF471: '樿' // U+6A3F <cjk>
	0xF472: '橆' // U+6A46 <cjk>
	0xF473: '橉' // U+6A49 <cjk>
	0xF474: '橺' // U+6A7A <cjk>
	0xF475: '橎' // U+6A4E <cjk>
	0xF476: '橒' // U+6A52 <cjk>
	0xF477: '橤' // U+6A64 <cjk>
	0xF478: '𣜌' // U+2370C <cjk>
	0xF479: '橾' // U+6A7E <cjk>
	0xF47A: '檃' // U+6A83 <cjk>
	0xF47B: '檋' // U+6A8B <cjk>
	0xF47C: '㯰' // U+3BF0 <cjk>
	0xF47D: '檑' // U+6A91 <cjk>
	0xF47E: '檟' // U+6A9F <cjk>
	0xF480: '檡' // U+6AA1 <cjk>
	0xF481: '𣝤' // U+23764 <cjk>
	0xF482: '檫' // U+6AAB <cjk>
	0xF483: '檽' // U+6ABD <cjk>
	0xF484: '櫆' // U+6AC6 <cjk>
	0xF485: '櫔' // U+6AD4 <cjk>
	0xF486: '櫐' // U+6AD0 <cjk>
	0xF487: '櫜' // U+6ADC <cjk>
	0xF488: '櫝' // U+6ADD <cjk>
	0xF489: '𣟿' // U+237FF <cjk>
	0xF48A: '𣟧' // U+237E7 <cjk>
	0xF48B: '櫬' // U+6AEC <cjk>
	0xF48C: '櫱' // U+6AF1 <cjk>
	0xF48D: '櫲' // U+6AF2 <cjk>
	0xF48E: '櫳' // U+6AF3 <cjk>
	0xF48F: '櫽' // U+6AFD <cjk>
	0xF490: '𣠤' // U+23824 <cjk>
	0xF491: '欋' // U+6B0B <cjk>
	0xF492: '欏' // U+6B0F <cjk>
	0xF493: '欐' // U+6B10 <cjk>
	0xF494: '欑' // U+6B11 <cjk>
	0xF495: '𣠽' // U+2383D <cjk>
	0xF496: '欗' // U+6B17 <cjk>
	0xF497: '㰦' // U+3C26 <cjk>
	0xF498: '欯' // U+6B2F <cjk>
	0xF499: '歊' // U+6B4A <cjk>
	0xF49A: '歘' // U+6B58 <cjk>
	0xF49B: '歬' // U+6B6C <cjk>
	0xF49C: '歵' // U+6B75 <cjk>
	0xF49D: '歺' // U+6B7A <cjk>
	0xF49E: '殁' // U+6B81 <cjk>
	0xF49F: '殛' // U+6B9B <cjk>
	0xF4A0: '殮' // U+6BAE <cjk>
	0xF4A1: '𣪘' // U+23A98 <cjk>
	0xF4A2: '殽' // U+6BBD <cjk>
	0xF4A3: '殾' // U+6BBE <cjk>
	0xF4A4: '毇' // U+6BC7 <cjk>
	0xF4A5: '毈' // U+6BC8 <cjk>
	0xF4A6: '毉' // U+6BC9 <cjk>
	0xF4A7: '毚' // U+6BDA <cjk>
	0xF4A8: '毦' // U+6BE6 <cjk>
	0xF4A9: '毧' // U+6BE7 <cjk>
	0xF4AA: '毮' // U+6BEE <cjk>
	0xF4AB: '毱' // U+6BF1 <cjk>
	0xF4AC: '氂' // U+6C02 <cjk>
	0xF4AD: '氊' // U+6C0A <cjk>
	0xF4AE: '氎' // U+6C0E <cjk>
	0xF4AF: '氵' // U+6C35 <cjk>
	0xF4B0: '氶' // U+6C36 <cjk>
	0xF4B1: '氺' // U+6C3A <cjk>
	0xF4B2: '𣱿' // U+23C7F <cjk>
	0xF4B3: '氿' // U+6C3F <cjk>
	0xF4B4: '汍' // U+6C4D <cjk>
	0xF4B5: '汛' // U+6C5B <cjk>
	0xF4B6: '汭' // U+6C6D <cjk>
	0xF4B7: '沄' // U+6C84 <cjk>
	0xF4B8: '沉' // U+6C89 <cjk>
	0xF4B9: '㳃' // U+3CC3 <cjk>
	0xF4BA: '沔' // U+6C94 <cjk>
	0xF4BB: '沕' // U+6C95 <cjk>
	0xF4BC: '沗' // U+6C97 <cjk>
	0xF4BD: '沭' // U+6CAD <cjk>
	0xF4BE: '泂' // U+6CC2 <cjk>
	0xF4BF: '泐' // U+6CD0 <cjk>
	0xF4C0: '㳒' // U+3CD2 <cjk>
	0xF4C1: '泖' // U+6CD6 <cjk>
	0xF4C2: '泚' // U+6CDA <cjk>
	0xF4C3: '泜' // U+6CDC <cjk>
	0xF4C4: '泩' // U+6CE9 <cjk>
	0xF4C5: '泬' // U+6CEC <cjk>
	0xF4C6: '泭' // U+6CED <cjk>
	0xF4C7: '𣴀' // U+23D00 <cjk>
	0xF4C8: '洀' // U+6D00 <cjk>
	0xF4C9: '洊' // U+6D0A <cjk>
	0xF4CA: '洤' // U+6D24 <cjk>
	0xF4CB: '洦' // U+6D26 <cjk>
	0xF4CC: '洧' // U+6D27 <cjk>
	0xF4CD: '汧' // U+6C67 <cjk>
	0xF4CE: '洯' // U+6D2F <cjk>
	0xF4CF: '洼' // U+6D3C <cjk>
	0xF4D0: '浛' // U+6D5B <cjk>
	0xF4D1: '浞' // U+6D5E <cjk>
	0xF4D2: '浠' // U+6D60 <cjk>
	0xF4D3: '浰' // U+6D70 <cjk>
	0xF4D4: '涀' // U+6D80 <cjk>
	0xF4D5: '涁' // U+6D81 <cjk>
	0xF4D6: '涊' // U+6D8A <cjk>
	0xF4D7: '涍' // U+6D8D <cjk>
	0xF4D8: '涑' // U+6D91 <cjk>
	0xF4D9: '涘' // U+6D98 <cjk>
	0xF4DA: '𣵀' // U+23D40 <cjk>
	0xF4DB: '渗' // U+6E17 <cjk>
	0xF4DC: '𣷺' // U+23DFA <cjk>
	0xF4DD: '𣷹' // U+23DF9 <cjk>
	0xF4DE: '𣷓' // U+23DD3 <cjk>
	0xF4DF: '涫' // U+6DAB <cjk>
	0xF4E0: '涮' // U+6DAE <cjk>
	0xF4E1: '涴' // U+6DB4 <cjk>
	0xF4E2: '淂' // U+6DC2 <cjk>
	0xF4E3: '洴' // U+6D34 <cjk>
	0xF4E4: '淈' // U+6DC8 <cjk>
	0xF4E5: '淎' // U+6DCE <cjk>
	0xF4E6: '淏' // U+6DCF <cjk>
	0xF4E7: '淐' // U+6DD0 <cjk>
	0xF4E8: '淟' // U+6DDF <cjk>
	0xF4E9: '淩' // U+6DE9 <cjk>
	0xF4EA: '淶' // U+6DF6 <cjk>
	0xF4EB: '渶' // U+6E36 <cjk>
	0xF4EC: '渞' // U+6E1E <cjk>
	0xF4ED: '渢' // U+6E22 <cjk>
	0xF4EE: '渧' // U+6E27 <cjk>
	0xF4EF: '㴑' // U+3D11 <cjk>
	0xF4F0: '渲' // U+6E32 <cjk>
	0xF4F1: '渼' // U+6E3C <cjk>
	0xF4F2: '湈' // U+6E48 <cjk>
	0xF4F3: '湉' // U+6E49 <cjk>
	0xF4F4: '湋' // U+6E4B <cjk>
	0xF4F5: '湌' // U+6E4C <cjk>
	0xF4F6: '湏' // U+6E4F <cjk>
	0xF4F7: '湑' // U+6E51 <cjk>
	0xF4F8: '湓' // U+6E53 <cjk>
	0xF4F9: '湔' // U+6E54 <cjk>
	0xF4FA: '湗' // U+6E57 <cjk>
	0xF4FB: '湣' // U+6E63 <cjk>
	0xF4FC: '㴞' // U+3D1E <cjk>
	0xF540: '溓' // U+6E93 <cjk>
	0xF541: '溧' // U+6EA7 <cjk>
	0xF542: '溴' // U+6EB4 <cjk>
	0xF543: '溿' // U+6EBF <cjk>
	0xF544: '滃' // U+6EC3 <cjk>
	0xF545: '滊' // U+6ECA <cjk>
	0xF546: '滙' // U+6ED9 <cjk>
	0xF547: '漵' // U+6F35 <cjk>
	0xF548: '滫' // U+6EEB <cjk>
	0xF549: '滹' // U+6EF9 <cjk>
	0xF54A: '滻' // U+6EFB <cjk>
	0xF54B: '漊' // U+6F0A <cjk>
	0xF54C: '漌' // U+6F0C <cjk>
	0xF54D: '漘' // U+6F18 <cjk>
	0xF54E: '漥' // U+6F25 <cjk>
	0xF54F: '漶' // U+6F36 <cjk>
	0xF550: '漼' // U+6F3C <cjk>
	0xF551: '𣽾' // U+23F7E <cjk>
	0xF552: '潒' // U+6F52 <cjk>
	0xF553: '潗' // U+6F57 <cjk>
	0xF554: '潚' // U+6F5A <cjk>
	0xF555: '潠' // U+6F60 <cjk>
	0xF556: '潨' // U+6F68 <cjk>
	0xF557: '澘' // U+6F98 <cjk>
	0xF558: '潽' // U+6F7D <cjk>
	0xF559: '澐' // U+6F90 <cjk>
	0xF55A: '澖' // U+6F96 <cjk>
	0xF55B: '澾' // U+6FBE <cjk>
	0xF55C: '澟' // U+6F9F <cjk>
	0xF55D: '澥' // U+6FA5 <cjk>
	0xF55E: '澯' // U+6FAF <cjk>
	0xF55F: '㵤' // U+3D64 <cjk>
	0xF560: '澵' // U+6FB5 <cjk>
	0xF561: '濈' // U+6FC8 <cjk>
	0xF562: '濉' // U+6FC9 <cjk>
	0xF563: '濚' // U+6FDA <cjk>
	0xF564: '濞' // U+6FDE <cjk>
	0xF565: '濩' // U+6FE9 <cjk>
	0xF566: '𤂖' // U+24096 <cjk>
	0xF567: '濼' // U+6FFC <cjk>
	0xF568: '瀀' // U+7000 <cjk>
	0xF569: '瀇' // U+7007 <cjk>
	0xF56A: '瀊' // U+700A <cjk>
	0xF56B: '瀣' // U+7023 <cjk>
	0xF56C: '𤄃' // U+24103 <cjk>
	0xF56D: '瀹' // U+7039 <cjk>
	0xF56E: '瀺' // U+703A <cjk>
	0xF56F: '瀼' // U+703C <cjk>
	0xF570: '灃' // U+7043 <cjk>
	0xF571: '灇' // U+7047 <cjk>
	0xF572: '灋' // U+704B <cjk>
	0xF573: '㶚' // U+3D9A <cjk>
	0xF574: '灔' // U+7054 <cjk>
	0xF575: '灥' // U+7065 <cjk>
	0xF576: '灩' // U+7069 <cjk>
	0xF577: '灬' // U+706C <cjk>
	0xF578: '灮' // U+706E <cjk>
	0xF579: '灶' // U+7076 <cjk>
	0xF57A: '灾' // U+707E <cjk>
	0xF57B: '炁' // U+7081 <cjk>
	0xF57C: '炆' // U+7086 <cjk>
	0xF57D: '炕' // U+7095 <cjk>
	0xF57E: '炗' // U+7097 <cjk>
	0xF580: '炻' // U+70BB <cjk>
	0xF581: '𤇆' // U+241C6 <cjk>
	0xF582: '炟' // U+709F <cjk>
	0xF583: '炱' // U+70B1 <cjk>
	0xF584: '𤇾' // U+241FE <cjk>
	0xF585: '烬' // U+70EC <cjk>
	0xF586: '烊' // U+70CA <cjk>
	0xF587: '烑' // U+70D1 <cjk>
	0xF588: '烓' // U+70D3 <cjk>
	0xF589: '烜' // U+70DC <cjk>
	0xF58A: '焃' // U+7103 <cjk>
	0xF58B: '焄' // U+7104 <cjk>
	0xF58C: '焆' // U+7106 <cjk>
	0xF58D: '焇' // U+7107 <cjk>
	0xF58E: '焈' // U+7108 <cjk>
	0xF58F: '焌' // U+710C <cjk>
	0xF590: '㷀' // U+3DC0 <cjk>
	0xF591: '焯' // U+712F <cjk>
	0xF592: '焱' // U+7131 <cjk>
	0xF593: '煐' // U+7150 <cjk>
	0xF594: '煊' // U+714A <cjk>
	0xF595: '煓' // U+7153 <cjk>
	0xF596: '煞' // U+715E <cjk>
	0xF597: '㷔' // U+3DD4 <cjk>
	0xF598: '熖' // U+7196 <cjk>
	0xF599: '熀' // U+7180 <cjk>
	0xF59A: '熛' // U+719B <cjk>
	0xF59B: '熠' // U+71A0 <cjk>
	0xF59C: '熢' // U+71A2 <cjk>
	0xF59D: '熮' // U+71AE <cjk>
	0xF59E: '熯' // U+71AF <cjk>
	0xF59F: '熳' // U+71B3 <cjk>
	0xF5A0: '𤎼' // U+243BC <cjk>
	0xF5A1: '燋' // U+71CB <cjk>
	0xF5A2: '燓' // U+71D3 <cjk>
	0xF5A3: '燙' // U+71D9 <cjk>
	0xF5A4: '燜' // U+71DC <cjk>
	0xF5A5: '爇' // U+7207 <cjk>
	0xF5A6: '㸅' // U+3E05 <cjk>
	0xF5A7: '爫' // U+FA49 CJK COMPATIBILITY IDEOGRAPH-FA49
	0xF5A8: '爫' // U+722B <cjk>
	0xF5A9: '爴' // U+7234 <cjk>
	0xF5AA: '爸' // U+7238 <cjk>
	0xF5AB: '爹' // U+7239 <cjk>
	0xF5AC: '丬' // U+4E2C <cjk>
	0xF5AD: '牂' // U+7242 <cjk>
	0xF5AE: '牓' // U+7253 <cjk>
	0xF5AF: '牗' // U+7257 <cjk>
	0xF5B0: '牣' // U+7263 <cjk>
	0xF5B1: '𤘩' // U+24629 <cjk>
	0xF5B2: '牮' // U+726E <cjk>
	0xF5B3: '牯' // U+726F <cjk>
	0xF5B4: '牸' // U+7278 <cjk>
	0xF5B5: '牿' // U+727F <cjk>
	0xF5B6: '犎' // U+728E <cjk>
	0xF5B7: '𤚥' // U+246A5 <cjk>
	0xF5B8: '犭' // U+72AD <cjk>
	0xF5B9: '犮' // U+72AE <cjk>
	0xF5BA: '犰' // U+72B0 <cjk>
	0xF5BB: '犱' // U+72B1 <cjk>
	0xF5BC: '狁' // U+72C1 <cjk>
	0xF5BD: '㹠' // U+3E60 <cjk>
	0xF5BE: '狌' // U+72CC <cjk>
	0xF5BF: '㹦' // U+3E66 <cjk>
	0xF5C0: '㹨' // U+3E68 <cjk>
	0xF5C1: '狳' // U+72F3 <cjk>
	0xF5C2: '狺' // U+72FA <cjk>
	0xF5C3: '猇' // U+7307 <cjk>
	0xF5C4: '猒' // U+7312 <cjk>
	0xF5C5: '猘' // U+7318 <cjk>
	0xF5C6: '猙' // U+7319 <cjk>
	0xF5C7: '㺃' // U+3E83 <cjk>
	0xF5C8: '猹' // U+7339 <cjk>
	0xF5C9: '猬' // U+732C <cjk>
	0xF5CA: '猱' // U+7331 <cjk>
	0xF5CB: '猳' // U+7333 <cjk>
	0xF5CC: '猽' // U+733D <cjk>
	0xF5CD: '獒' // U+7352 <cjk>
	0xF5CE: '㺔' // U+3E94 <cjk>
	0xF5CF: '獫' // U+736B <cjk>
	0xF5D0: '獬' // U+736C <cjk>
	0xF5D1: '𤢖' // U+24896 <cjk>
	0xF5D2: '獮' // U+736E <cjk>
	0xF5D3: '獯' // U+736F <cjk>
	0xF5D4: '獱' // U+7371 <cjk>
	0xF5D5: '獷' // U+7377 <cjk>
	0xF5D6: '玁' // U+7381 <cjk>
	0xF5D7: '玅' // U+7385 <cjk>
	0xF5D8: '玊' // U+738A <cjk>
	0xF5D9: '玔' // U+7394 <cjk>
	0xF5DA: '玘' // U+7398 <cjk>
	0xF5DB: '玜' // U+739C <cjk>
	0xF5DC: '玞' // U+739E <cjk>
	0xF5DD: '玥' // U+73A5 <cjk>
	0xF5DE: '玨' // U+73A8 <cjk>
	0xF5DF: '玵' // U+73B5 <cjk>
	0xF5E0: '玷' // U+73B7 <cjk>
	0xF5E1: '玹' // U+73B9 <cjk>
	0xF5E2: '玼' // U+73BC <cjk>
	0xF5E3: '玿' // U+73BF <cjk>
	0xF5E4: '珅' // U+73C5 <cjk>
	0xF5E5: '珋' // U+73CB <cjk>
	0xF5E6: '珡' // U+73E1 <cjk>
	0xF5E7: '珧' // U+73E7 <cjk>
	0xF5E8: '珹' // U+73F9 <cjk>
	0xF5E9: '琓' // U+7413 <cjk>
	0xF5EA: '珺' // U+73FA <cjk>
	0xF5EB: '琁' // U+7401 <cjk>
	0xF5EC: '琤' // U+7424 <cjk>
	0xF5ED: '琱' // U+7431 <cjk>
	0xF5EE: '琹' // U+7439 <cjk>
	0xF5EF: '瑓' // U+7453 <cjk>
	0xF5F0: '瑀' // U+7440 <cjk>
	0xF5F1: '瑃' // U+7443 <cjk>
	0xF5F2: '瑍' // U+744D <cjk>
	0xF5F3: '瑒' // U+7452 <cjk>
	0xF5F4: '瑝' // U+745D <cjk>
	0xF5F5: '瑱' // U+7471 <cjk>
	0xF5F6: '璁' // U+7481 <cjk>
	0xF5F7: '璅' // U+7485 <cjk>
	0xF5F8: '璈' // U+7488 <cjk>
	0xF5F9: '𤩍' // U+24A4D <cjk>
	0xF5FA: '璒' // U+7492 <cjk>
	0xF5FB: '璗' // U+7497 <cjk>
	0xF5FC: '璙' // U+7499 <cjk>
	0xF640: '璠' // U+74A0 <cjk>
	0xF641: '璡' // U+74A1 <cjk>
	0xF642: '璥' // U+74A5 <cjk>
	0xF643: '璪' // U+74AA <cjk>
	0xF644: '璫' // U+74AB <cjk>
	0xF645: '璹' // U+74B9 <cjk>
	0xF646: '璻' // U+74BB <cjk>
	0xF647: '璺' // U+74BA <cjk>
	0xF648: '瓖' // U+74D6 <cjk>
	0xF649: '瓘' // U+74D8 <cjk>
	0xF64A: '瓞' // U+74DE <cjk>
	0xF64B: '瓯' // U+74EF <cjk>
	0xF64C: '瓫' // U+74EB <cjk>
	0xF64D: '𤭖' // U+24B56 <cjk>
	0xF64E: '瓺' // U+74FA <cjk>
	0xF64F: '𤭯' // U+24B6F <cjk>
	0xF650: '甠' // U+7520 <cjk>
	0xF651: '甤' // U+7524 <cjk>
	0xF652: '甪' // U+752A <cjk>
	0xF653: '㽗' // U+3F57 <cjk>
	0xF654: '𤰖' // U+24C16 <cjk>
	0xF655: '甽' // U+753D <cjk>
	0xF656: '甾' // U+753E <cjk>
	0xF657: '畀' // U+7540 <cjk>
	0xF658: '畈' // U+7548 <cjk>
	0xF659: '畎' // U+754E <cjk>
	0xF65A: '畐' // U+7550 <cjk>
	0xF65B: '畒' // U+7552 <cjk>
	0xF65C: '畬' // U+756C <cjk>
	0xF65D: '畲' // U+7572 <cjk>
	0xF65E: '畱' // U+7571 <cjk>
	0xF65F: '畺' // U+757A <cjk>
	0xF660: '畽' // U+757D <cjk>
	0xF661: '畾' // U+757E <cjk>
	0xF662: '疁' // U+7581 <cjk>
	0xF663: '𤴔' // U+24D14 <cjk>
	0xF664: '疌' // U+758C <cjk>
	0xF665: '㽵' // U+3F75 <cjk>
	0xF666: '疢' // U+75A2 <cjk>
	0xF667: '㽷' // U+3F77 <cjk>
	0xF668: '疰' // U+75B0 <cjk>
	0xF669: '疷' // U+75B7 <cjk>
	0xF66A: '疿' // U+75BF <cjk>
	0xF66B: '痀' // U+75C0 <cjk>
	0xF66C: '痆' // U+75C6 <cjk>
	0xF66D: '痏' // U+75CF <cjk>
	0xF66E: '痓' // U+75D3 <cjk>
	0xF66F: '痝' // U+75DD <cjk>
	0xF670: '痟' // U+75DF <cjk>
	0xF671: '痠' // U+75E0 <cjk>
	0xF672: '痧' // U+75E7 <cjk>
	0xF673: '痬' // U+75EC <cjk>
	0xF674: '痮' // U+75EE <cjk>
	0xF675: '痱' // U+75F1 <cjk>
	0xF676: '痹' // U+75F9 <cjk>
	0xF677: '瘃' // U+7603 <cjk>
	0xF678: '瘘' // U+7618 <cjk>
	0xF679: '瘇' // U+7607 <cjk>
	0xF67A: '瘏' // U+760F <cjk>
	0xF67B: '㾮' // U+3FAE <cjk>
	0xF67C: '𤸎' // U+24E0E <cjk>
	0xF67D: '瘓' // U+7613 <cjk>
	0xF67E: '瘛' // U+761B <cjk>
	0xF680: '瘜' // U+761C <cjk>
	0xF681: '𤸷' // U+24E37 <cjk>
	0xF682: '瘥' // U+7625 <cjk>
	0xF683: '瘨' // U+7628 <cjk>
	0xF684: '瘼' // U+763C <cjk>
	0xF685: '瘳' // U+7633 <cjk>
	0xF686: '𤹪' // U+24E6A <cjk>
	0xF687: '㿉' // U+3FC9 <cjk>
	0xF688: '癁' // U+7641 <cjk>
	0xF689: '𤺋' // U+24E8B <cjk>
	0xF68A: '癉' // U+7649 <cjk>
	0xF68B: '癕' // U+7655 <cjk>
	0xF68C: '㿗' // U+3FD7 <cjk>
	0xF68D: '癮' // U+766E <cjk>
	0xF68E: '皕' // U+7695 <cjk>
	0xF68F: '皜' // U+769C <cjk>
	0xF690: '皡' // U+76A1 <cjk>
	0xF691: '皠' // U+76A0 <cjk>
	0xF692: '皧' // U+76A7 <cjk>
	0xF693: '皨' // U+76A8 <cjk>
	0xF694: '皯' // U+76AF <cjk>
	0xF695: '𥁊' // U+2504A <cjk>
	0xF696: '盉' // U+76C9 <cjk>
	0xF697: '𥁕' // U+25055 <cjk>
	0xF698: '盨' // U+76E8 <cjk>
	0xF699: '盬' // U+76EC <cjk>
	0xF69A: '𥄢' // U+25122 <cjk>
	0xF69B: '眗' // U+7717 <cjk>
	0xF69C: '眚' // U+771A <cjk>
	0xF69D: '眭' // U+772D <cjk>
	0xF69E: '眵' // U+7735 <cjk>
	0xF69F: '𥆩' // U+251A9 <cjk>
	0xF6A0: '䀹' // U+4039 <cjk>
	0xF6A1: '𥇥' // U+251E5 <cjk>
	0xF6A2: '𥇍' // U+251CD <cjk>
	0xF6A3: '睘' // U+7758 <cjk>
	0xF6A4: '睠' // U+7760 <cjk>
	0xF6A5: '睪' // U+776A <cjk>
	0xF6A6: '𥈞' // U+2521E <cjk>
	0xF6A7: '睲' // U+7772 <cjk>
	0xF6A8: '睼' // U+777C <cjk>
	0xF6A9: '睽' // U+777D <cjk>
	0xF6AA: '𥉌' // U+2524C <cjk>
	0xF6AB: '䁘' // U+4058 <cjk>
	0xF6AC: '瞚' // U+779A <cjk>
	0xF6AD: '瞟' // U+779F <cjk>
	0xF6AE: '瞢' // U+77A2 <cjk>
	0xF6AF: '瞤' // U+77A4 <cjk>
	0xF6B0: '瞩' // U+77A9 <cjk>
	0xF6B1: '矞' // U+77DE <cjk>
	0xF6B2: '矟' // U+77DF <cjk>
	0xF6B3: '矤' // U+77E4 <cjk>
	0xF6B4: '矦' // U+77E6 <cjk>
	0xF6B5: '矪' // U+77EA <cjk>
	0xF6B6: '矬' // U+77EC <cjk>
	0xF6B7: '䂓' // U+4093 <cjk>
	0xF6B8: '矰' // U+77F0 <cjk>
	0xF6B9: '矴' // U+77F4 <cjk>
	0xF6BA: '矻' // U+77FB <cjk>
	0xF6BB: '𥐮' // U+2542E <cjk>
	0xF6BC: '砅' // U+7805 <cjk>
	0xF6BD: '砆' // U+7806 <cjk>
	0xF6BE: '砉' // U+7809 <cjk>
	0xF6BF: '砍' // U+780D <cjk>
	0xF6C0: '砙' // U+7819 <cjk>
	0xF6C1: '砡' // U+7821 <cjk>
	0xF6C2: '砬' // U+782C <cjk>
	0xF6C3: '硇' // U+7847 <cjk>
	0xF6C4: '硤' // U+7864 <cjk>
	0xF6C5: '硪' // U+786A <cjk>
	0xF6C6: '𥓙' // U+254D9 <cjk>
	0xF6C7: '碊' // U+788A <cjk>
	0xF6C8: '碔' // U+7894 <cjk>
	0xF6C9: '碤' // U+78A4 <cjk>
	0xF6CA: '碝' // U+789D <cjk>
	0xF6CB: '碞' // U+789E <cjk>
	0xF6CC: '碟' // U+789F <cjk>
	0xF6CD: '碻' // U+78BB <cjk>
	0xF6CE: '磈' // U+78C8 <cjk>
	0xF6CF: '磌' // U+78CC <cjk>
	0xF6D0: '磎' // U+78CE <cjk>
	0xF6D1: '磕' // U+78D5 <cjk>
	0xF6D2: '磠' // U+78E0 <cjk>
	0xF6D3: '磡' // U+78E1 <cjk>
	0xF6D4: '磦' // U+78E6 <cjk>
	0xF6D5: '磹' // U+78F9 <cjk>
	0xF6D6: '磺' // U+78FA <cjk>
	0xF6D7: '磻' // U+78FB <cjk>
	0xF6D8: '磾' // U+78FE <cjk>
	0xF6D9: '𥖧' // U+255A7 <cjk>
	0xF6DA: '礐' // U+7910 <cjk>
	0xF6DB: '礛' // U+791B <cjk>
	0xF6DC: '礰' // U+7930 <cjk>
	0xF6DD: '礥' // U+7925 <cjk>
	0xF6DE: '礻' // U+793B <cjk>
	0xF6DF: '祊' // U+794A <cjk>
	0xF6E0: '祘' // U+7958 <cjk>
	0xF6E1: '祛' // U+795B <cjk>
	0xF6E2: '䄅' // U+4105 <cjk>
	0xF6E3: '祧' // U+7967 <cjk>
	0xF6E4: '祲' // U+7972 <cjk>
	0xF6E5: '禔' // U+7994 <cjk>
	0xF6E6: '禕' // U+7995 <cjk>
	0xF6E7: '禖' // U+7996 <cjk>
	0xF6E8: '禛' // U+799B <cjk>
	0xF6E9: '禡' // U+79A1 <cjk>
	0xF6EA: '禩' // U+79A9 <cjk>
	0xF6EB: '禴' // U+79B4 <cjk>
	0xF6EC: '离' // U+79BB <cjk>
	0xF6ED: '秂' // U+79C2 <cjk>
	0xF6EE: '秇' // U+79C7 <cjk>
	0xF6EF: '秌' // U+79CC <cjk>
	0xF6F0: '种' // U+79CD <cjk>
	0xF6F1: '秖' // U+79D6 <cjk>
	0xF6F2: '䅈' // U+4148 <cjk>
	0xF6F3: '𥞩' // U+257A9 <cjk>
	0xF6F4: '𥞴' // U+257B4 <cjk>
	0xF6F5: '䅏' // U+414F <cjk>
	0xF6F6: '稊' // U+7A0A <cjk>
	0xF6F7: '稑' // U+7A11 <cjk>
	0xF6F8: '稕' // U+7A15 <cjk>
	0xF6F9: '稛' // U+7A1B <cjk>
	0xF6FA: '稞' // U+7A1E <cjk>
	0xF6FB: '䅣' // U+4163 <cjk>
	0xF6FC: '稭' // U+7A2D <cjk>
	0xF740: '稸' // U+7A38 <cjk>
	0xF741: '穇' // U+7A47 <cjk>
	0xF742: '穌' // U+7A4C <cjk>
	0xF743: '穖' // U+7A56 <cjk>
	0xF744: '穙' // U+7A59 <cjk>
	0xF745: '穜' // U+7A5C <cjk>
	0xF746: '穟' // U+7A5F <cjk>
	0xF747: '穠' // U+7A60 <cjk>
	0xF748: '穧' // U+7A67 <cjk>
	0xF749: '穪' // U+7A6A <cjk>
	0xF74A: '穵' // U+7A75 <cjk>
	0xF74B: '穸' // U+7A78 <cjk>
	0xF74C: '窂' // U+7A82 <cjk>
	0xF74D: '窊' // U+7A8A <cjk>
	0xF74E: '窐' // U+7A90 <cjk>
	0xF74F: '窣' // U+7AA3 <cjk>
	0xF750: '窬' // U+7AAC <cjk>
	0xF751: '𥧔' // U+259D4 <cjk>
	0xF752: '䆴' // U+41B4 <cjk>
	0xF753: '窹' // U+7AB9 <cjk>
	0xF754: '窼' // U+7ABC <cjk>
	0xF755: '窾' // U+7ABE <cjk>
	0xF756: '䆿' // U+41BF <cjk>
	0xF757: '竌' // U+7ACC <cjk>
	0xF758: '竑' // U+7AD1 <cjk>
	0xF759: '竧' // U+7AE7 <cjk>
	0xF75A: '竨' // U+7AE8 <cjk>
	0xF75B: '竴' // U+7AF4 <cjk>
	0xF75C: '𥫤' // U+25AE4 <cjk>
	0xF75D: '𥫣' // U+25AE3 <cjk>
	0xF75E: '笇' // U+7B07 <cjk>
	0xF75F: '𥫱' // U+25AF1 <cjk>
	0xF760: '笽' // U+7B3D <cjk>
	0xF761: '笧' // U+7B27 <cjk>
	0xF762: '笪' // U+7B2A <cjk>
	0xF763: '笮' // U+7B2E <cjk>
	0xF764: '笯' // U+7B2F <cjk>
	0xF765: '笱' // U+7B31 <cjk>
	0xF766: '䇦' // U+41E6 <cjk>
	0xF767: '䇳' // U+41F3 <cjk>
	0xF768: '筿' // U+7B7F <cjk>
	0xF769: '筁' // U+7B41 <cjk>
	0xF76A: '䇮' // U+41EE <cjk>
	0xF76B: '筕' // U+7B55 <cjk>
	0xF76C: '筹' // U+7B79 <cjk>
	0xF76D: '筤' // U+7B64 <cjk>
	0xF76E: '筦' // U+7B66 <cjk>
	0xF76F: '筩' // U+7B69 <cjk>
	0xF770: '筳' // U+7B73 <cjk>
	0xF771: '𥮲' // U+25BB2 <cjk>
	0xF772: '䈇' // U+4207 <cjk>
	0xF773: '箐' // U+7B90 <cjk>
	0xF774: '箑' // U+7B91 <cjk>
	0xF775: '箛' // U+7B9B <cjk>
	0xF776: '䈎' // U+420E <cjk>
	0xF777: '箯' // U+7BAF <cjk>
	0xF778: '箵' // U+7BB5 <cjk>
	0xF779: '箼' // U+7BBC <cjk>
	0xF77A: '篅' // U+7BC5 <cjk>
	0xF77B: '篊' // U+7BCA <cjk>
	0xF77C: '𥱋' // U+25C4B <cjk>
	0xF77D: '𥱤' // U+25C64 <cjk>
	0xF77E: '篔' // U+7BD4 <cjk>
	0xF780: '篖' // U+7BD6 <cjk>
	0xF781: '篚' // U+7BDA <cjk>
	0xF782: '篪' // U+7BEA <cjk>
	0xF783: '篰' // U+7BF0 <cjk>
	0xF784: '簃' // U+7C03 <cjk>
	0xF785: '簋' // U+7C0B <cjk>
	0xF786: '簎' // U+7C0E <cjk>
	0xF787: '簏' // U+7C0F <cjk>
	0xF788: '簦' // U+7C26 <cjk>
	0xF789: '籅' // U+7C45 <cjk>
	0xF78A: '籊' // U+7C4A <cjk>
	0xF78B: '籑' // U+7C51 <cjk>
	0xF78C: '籗' // U+7C57 <cjk>
	0xF78D: '籞' // U+7C5E <cjk>
	0xF78E: '籡' // U+7C61 <cjk>
	0xF78F: '籩' // U+7C69 <cjk>
	0xF790: '籮' // U+7C6E <cjk>
	0xF791: '籯' // U+7C6F <cjk>
	0xF792: '籰' // U+7C70 <cjk>
	0xF793: '𥸮' // U+25E2E <cjk>
	0xF794: '𥹖' // U+25E56 <cjk>
	0xF795: '𥹥' // U+25E65 <cjk>
	0xF796: '粦' // U+7CA6 <cjk>
	0xF797: '𥹢' // U+25E62 <cjk>
	0xF798: '粶' // U+7CB6 <cjk>
	0xF799: '粷' // U+7CB7 <cjk>
	0xF79A: '粿' // U+7CBF <cjk>
	0xF79B: '𥻘' // U+25ED8 <cjk>
	0xF79C: '糄' // U+7CC4 <cjk>
	0xF79D: '𥻂' // U+25EC2 <cjk>
	0xF79E: '糈' // U+7CC8 <cjk>
	0xF79F: '糍' // U+7CCD <cjk>
	0xF7A0: '𥻨' // U+25EE8 <cjk>
	0xF7A1: '糗' // U+7CD7 <cjk>
	0xF7A2: '𥼣' // U+25F23 <cjk>
	0xF7A3: '糦' // U+7CE6 <cjk>
	0xF7A4: '糫' // U+7CEB <cjk>
	0xF7A5: '𥽜' // U+25F5C <cjk>
	0xF7A6: '糵' // U+7CF5 <cjk>
	0xF7A7: '紃' // U+7D03 <cjk>
	0xF7A8: '紉' // U+7D09 <cjk>
	0xF7A9: '䋆' // U+42C6 <cjk>
	0xF7AA: '紒' // U+7D12 <cjk>
	0xF7AB: '紞' // U+7D1E <cjk>
	0xF7AC: '𥿠' // U+25FE0 <cjk>
	0xF7AD: '𥿔' // U+25FD4 <cjk>
	0xF7AE: '紽' // U+7D3D <cjk>
	0xF7AF: '紾' // U+7D3E <cjk>
	0xF7B0: '絀' // U+7D40 <cjk>
	0xF7B1: '絇' // U+7D47 <cjk>
	0xF7B2: '𦀌' // U+2600C <cjk>
	0xF7B3: '𥿻' // U+25FFB <cjk>
	0xF7B4: '䋖' // U+42D6 <cjk>
	0xF7B5: '絙' // U+7D59 <cjk>
	0xF7B6: '絚' // U+7D5A <cjk>
	0xF7B7: '絪' // U+7D6A <cjk>
	0xF7B8: '絰' // U+7D70 <cjk>
	0xF7B9: '䋝' // U+42DD <cjk>
	0xF7BA: '絿' // U+7D7F <cjk>
	0xF7BB: '𦀗' // U+26017 <cjk>
	0xF7BC: '綆' // U+7D86 <cjk>
	0xF7BD: '綈' // U+7D88 <cjk>
	0xF7BE: '綌' // U+7D8C <cjk>
	0xF7BF: '綗' // U+7D97 <cjk>
	0xF7C0: '𦁠' // U+26060 <cjk>
	0xF7C1: '綝' // U+7D9D <cjk>
	0xF7C2: '綧' // U+7DA7 <cjk>
	0xF7C3: '綪' // U+7DAA <cjk>
	0xF7C4: '綶' // U+7DB6 <cjk>
	0xF7C5: '綷' // U+7DB7 <cjk>
	0xF7C6: '緀' // U+7DC0 <cjk>
	0xF7C7: '緗' // U+7DD7 <cjk>
	0xF7C8: '緙' // U+7DD9 <cjk>
	0xF7C9: '緦' // U+7DE6 <cjk>
	0xF7CA: '緱' // U+7DF1 <cjk>
	0xF7CB: '緹' // U+7DF9 <cjk>
	0xF7CC: '䌂' // U+4302 <cjk>
	0xF7CD: '𦃭' // U+260ED <cjk>
	0xF7CE: '縉' // U+FA58 CJK COMPATIBILITY IDEOGRAPH-FA58
	0xF7CF: '縐' // U+7E10 <cjk>
	0xF7D0: '縗' // U+7E17 <cjk>
	0xF7D1: '縝' // U+7E1D <cjk>
	0xF7D2: '縠' // U+7E20 <cjk>
	0xF7D3: '縧' // U+7E27 <cjk>
	0xF7D4: '縬' // U+7E2C <cjk>
	0xF7D5: '繅' // U+7E45 <cjk>
	0xF7D6: '繳' // U+7E73 <cjk>
	0xF7D7: '繵' // U+7E75 <cjk>
	0xF7D8: '繾' // U+7E7E <cjk>
	0xF7D9: '纆' // U+7E86 <cjk>
	0xF7DA: '纇' // U+7E87 <cjk>
	0xF7DB: '䌫' // U+432B <cjk>
	0xF7DC: '纑' // U+7E91 <cjk>
	0xF7DD: '纘' // U+7E98 <cjk>
	0xF7DE: '纚' // U+7E9A <cjk>
	0xF7DF: '䍃' // U+4343 <cjk>
	0xF7E0: '缼' // U+7F3C <cjk>
	0xF7E1: '缻' // U+7F3B <cjk>
	0xF7E2: '缾' // U+7F3E <cjk>
	0xF7E3: '罃' // U+7F43 <cjk>
	0xF7E4: '罄' // U+7F44 <cjk>
	0xF7E5: '罏' // U+7F4F <cjk>
	0xF7E6: '㓁' // U+34C1 <cjk>
	0xF7E7: '𦉰' // U+26270 <cjk>
	0xF7E8: '罒' // U+7F52 <cjk>
	0xF7E9: '𦊆' // U+26286 <cjk>
	0xF7EA: '罡' // U+7F61 <cjk>
	0xF7EB: '罣' // U+7F63 <cjk>
	0xF7EC: '罤' // U+7F64 <cjk>
	0xF7ED: '罭' // U+7F6D <cjk>
	0xF7EE: '罽' // U+7F7D <cjk>
	0xF7EF: '罾' // U+7F7E <cjk>
	0xF7F0: '𦍌' // U+2634C <cjk>
	0xF7F1: '羐' // U+7F90 <cjk>
	0xF7F2: '养' // U+517B <cjk>
	0xF7F3: '𣴎' // U+23D0E <cjk>
	0xF7F4: '羖' // U+7F96 <cjk>
	0xF7F5: '羜' // U+7F9C <cjk>
	0xF7F6: '羭' // U+7FAD <cjk>
	0xF7F7: '𦐂' // U+26402 <cjk>
	0xF7F8: '翃' // U+7FC3 <cjk>
	0xF7F9: '翏' // U+7FCF <cjk>
	0xF7FA: '翣' // U+7FE3 <cjk>
	0xF7FB: '翥' // U+7FE5 <cjk>
	0xF7FC: '翯' // U+7FEF <cjk>
	0xF840: '翲' // U+7FF2 <cjk>
	0xF841: '耂' // U+8002 <cjk>
	0xF842: '耊' // U+800A <cjk>
	0xF843: '耈' // U+8008 <cjk>
	0xF844: '耎' // U+800E <cjk>
	0xF845: '耑' // U+8011 <cjk>
	0xF846: '耖' // U+8016 <cjk>
	0xF847: '耤' // U+8024 <cjk>
	0xF848: '耬' // U+802C <cjk>
	0xF849: '耰' // U+8030 <cjk>
	0xF84A: '聃' // U+8043 <cjk>
	0xF84B: '聦' // U+8066 <cjk>
	0xF84C: '聱' // U+8071 <cjk>
	0xF84D: '聵' // U+8075 <cjk>
	0xF84E: '聻' // U+807B <cjk>
	0xF84F: '肙' // U+8099 <cjk>
	0xF850: '肜' // U+809C <cjk>
	0xF851: '肤' // U+80A4 <cjk>
	0xF852: '肧' // U+80A7 <cjk>
	0xF853: '肸' // U+80B8 <cjk>
	0xF854: '𦙾' // U+2667E <cjk>
	0xF855: '胅' // U+80C5 <cjk>
	0xF856: '胕' // U+80D5 <cjk>
	0xF857: '胘' // U+80D8 <cjk>
	0xF858: '胦' // U+80E6 <cjk>
	0xF859: '𦚰' // U+266B0 <cjk>
	0xF85A: '脍' // U+810D <cjk>
	0xF85B: '胵' // U+80F5 <cjk>
	0xF85C: '胻' // U+80FB <cjk>
	0xF85D: '䏮' // U+43EE <cjk>
	0xF85E: '脵' // U+8135 <cjk>
	0xF85F: '脖' // U+8116 <cjk>
	0xF860: '脞' // U+811E <cjk>
	0xF861: '䏰' // U+43F0 <cjk>
	0xF862: '脤' // U+8124 <cjk>
	0xF863: '脧' // U+8127 <cjk>
	0xF864: '脬' // U+812C <cjk>
	0xF865: '𦜝' // U+2671D <cjk>
	0xF866: '脽' // U+813D <cjk>
	0xF867: '䐈' // U+4408 <cjk>
	0xF868: '腩' // U+8169 <cjk>
	0xF869: '䐗' // U+4417 <cjk>
	0xF86A: '膁' // U+8181 <cjk>
	0xF86B: '䐜' // U+441C <cjk>
	0xF86C: '膄' // U+8184 <cjk>
	0xF86D: '膅' // U+8185 <cjk>
	0xF86E: '䐢' // U+4422 <cjk>
	0xF86F: '膘' // U+8198 <cjk>
	0xF870: '膲' // U+81B2 <cjk>
	0xF871: '臁' // U+81C1 <cjk>
	0xF872: '臃' // U+81C3 <cjk>
	0xF873: '臖' // U+81D6 <cjk>
	0xF874: '臛' // U+81DB <cjk>
	0xF875: '𦣝' // U+268DD <cjk>
	0xF876: '臤' // U+81E4 <cjk>
	0xF877: '𦣪' // U+268EA <cjk>
	0xF878: '臬' // U+81EC <cjk>
	0xF879: '𦥑' // U+26951 <cjk>
	0xF87A: '臽' // U+81FD <cjk>
	0xF87B: '臿' // U+81FF <cjk>
	0xF87C: '𦥯' // U+2696F <cjk>
	0xF87D: '舄' // U+8204 <cjk>
	0xF87E: '𦧝' // U+269DD <cjk>
	0xF880: '舙' // U+8219 <cjk>
	0xF881: '舡' // U+8221 <cjk>
	0xF882: '舢' // U+8222 <cjk>
	0xF883: '𦨞' // U+26A1E <cjk>
	0xF884: '舲' // U+8232 <cjk>
	0xF885: '舴' // U+8234 <cjk>
	0xF886: '舼' // U+823C <cjk>
	0xF887: '艆' // U+8246 <cjk>
	0xF888: '艉' // U+8249 <cjk>
	0xF889: '艅' // U+8245 <cjk>
	0xF88A: '𦩘' // U+26A58 <cjk>
	0xF88B: '艋' // U+824B <cjk>
	0xF88C: '䑶' // U+4476 <cjk>
	0xF88D: '艏' // U+824F <cjk>
	0xF88E: '䑺' // U+447A <cjk>
	0xF88F: '艗' // U+8257 <cjk>
	0xF890: '𦪌' // U+26A8C <cjk>
	0xF891: '艜' // U+825C <cjk>
	0xF892: '艣' // U+8263 <cjk>
	0xF893: '𦪷' // U+26AB7 <cjk>
	0xF894: '艹' // U+FA5D CJK COMPATIBILITY IDEOGRAPH-FA5D
	0xF895: '艹' // U+FA5E CJK COMPATIBILITY IDEOGRAPH-FA5E
	0xF896: '艹' // U+8279 <cjk>
	0xF897: '䒑' // U+4491 <cjk>
	0xF898: '艽' // U+827D <cjk>
	0xF899: '艿' // U+827F <cjk>
	0xF89A: '芃' // U+8283 <cjk>
	0xF89B: '芊' // U+828A <cjk>
	0xF89C: '芓' // U+8293 <cjk>
	0xF89D: '芧' // U+82A7 <cjk>
	0xF89E: '芨' // U+82A8 <cjk>
	0xF89F: '芲' // U+82B2 <cjk>
	0xF8A0: '芴' // U+82B4 <cjk>
	0xF8A1: '芺' // U+82BA <cjk>
	0xF8A2: '芼' // U+82BC <cjk>
	0xF8A3: '苢' // U+82E2 <cjk>
	0xF8A4: '苨' // U+82E8 <cjk>
	0xF8A5: '苷' // U+82F7 <cjk>
	0xF8A6: '茇' // U+8307 <cjk>
	0xF8A7: '茈' // U+8308 <cjk>
	0xF8A8: '茌' // U+830C <cjk>
	0xF8A9: '荔' // U+8354 <cjk>
	0xF8AA: '茛' // U+831B <cjk>
	0xF8AB: '茝' // U+831D <cjk>
	0xF8AC: '茰' // U+8330 <cjk>
	0xF8AD: '茼' // U+833C <cjk>
	0xF8AE: '荄' // U+8344 <cjk>
	0xF8AF: '荗' // U+8357 <cjk>
	0xF8B0: '䒾' // U+44BE <cjk>
	0xF8B1: '荿' // U+837F <cjk>
	0xF8B2: '䓔' // U+44D4 <cjk>
	0xF8B3: '䒳' // U+44B3 <cjk>
	0xF8B4: '莍' // U+838D <cjk>
	0xF8B5: '莔' // U+8394 <cjk>
	0xF8B6: '莕' // U+8395 <cjk>
	0xF8B7: '莛' // U+839B <cjk>
	0xF8B8: '莝' // U+839D <cjk>
	0xF8B9: '菉' // U+83C9 <cjk>
	0xF8BA: '菐' // U+83D0 <cjk>
	0xF8BB: '菔' // U+83D4 <cjk>
	0xF8BC: '菝' // U+83DD <cjk>
	0xF8BD: '菥' // U+83E5 <cjk>
	0xF8BE: '菹' // U+83F9 <cjk>
	0xF8BF: '萏' // U+840F <cjk>
	0xF8C0: '萑' // U+8411 <cjk>
	0xF8C1: '萕' // U+8415 <cjk>
	0xF8C2: '𦱳' // U+26C73 <cjk>
	0xF8C3: '萗' // U+8417 <cjk>
	0xF8C4: '萹' // U+8439 <cjk>
	0xF8C5: '葊' // U+844A <cjk>
	0xF8C6: '葏' // U+844F <cjk>
	0xF8C7: '葑' // U+8451 <cjk>
	0xF8C8: '葒' // U+8452 <cjk>
	0xF8C9: '葙' // U+8459 <cjk>
	0xF8CA: '葚' // U+845A <cjk>
	0xF8CB: '葜' // U+845C <cjk>
	0xF8CC: '𦳝' // U+26CDD <cjk>
	0xF8CD: '葥' // U+8465 <cjk>
	0xF8CE: '葶' // U+8476 <cjk>
	0xF8CF: '葸' // U+8478 <cjk>
	0xF8D0: '葼' // U+847C <cjk>
	0xF8D1: '蒁' // U+8481 <cjk>
	0xF8D2: '䔍' // U+450D <cjk>
	0xF8D3: '蓜' // U+84DC <cjk>
	0xF8D4: '蒗' // U+8497 <cjk>
	0xF8D5: '蒦' // U+84A6 <cjk>
	0xF8D6: '蒾' // U+84BE <cjk>
	0xF8D7: '䔈' // U+4508 <cjk>
	0xF8D8: '蓎' // U+84CE <cjk>
	0xF8D9: '蓏' // U+84CF <cjk>
	0xF8DA: '蓓' // U+84D3 <cjk>
	0xF8DB: '𦹥' // U+26E65 <cjk>
	0xF8DC: '蓧' // U+84E7 <cjk>
	0xF8DD: '蓪' // U+84EA <cjk>
	0xF8DE: '蓯' // U+84EF <cjk>
	0xF8DF: '蓰' // U+84F0 <cjk>
	0xF8E0: '蓱' // U+84F1 <cjk>
	0xF8E1: '蓺' // U+84FA <cjk>
	0xF8E2: '蓽' // U+84FD <cjk>
	0xF8E3: '蔌' // U+850C <cjk>
	0xF8E4: '蔛' // U+851B <cjk>
	0xF8E5: '蔤' // U+8524 <cjk>
	0xF8E6: '蔥' // U+8525 <cjk>
	0xF8E7: '蔫' // U+852B <cjk>
	0xF8E8: '蔴' // U+8534 <cjk>
	0xF8E9: '蕏' // U+854F <cjk>
	0xF8EA: '蕯' // U+856F <cjk>
	0xF8EB: '䔥' // U+4525 <cjk>
	0xF8EC: '䕃' // U+4543 <cjk>
	0xF8ED: '蔾' // U+853E <cjk>
	0xF8EE: '蕑' // U+8551 <cjk>
	0xF8EF: '蕓' // U+8553 <cjk>
	0xF8F0: '蕞' // U+855E <cjk>
	0xF8F1: '蕡' // U+8561 <cjk>
	0xF8F2: '蕢' // U+8562 <cjk>
	0xF8F3: '𦾔' // U+26F94 <cjk>
	0xF8F4: '蕻' // U+857B <cjk>
	0xF8F5: '蕽' // U+857D <cjk>
	0xF8F6: '蕿' // U+857F <cjk>
	0xF8F7: '薁' // U+8581 <cjk>
	0xF8F8: '薆' // U+8586 <cjk>
	0xF8F9: '薓' // U+8593 <cjk>
	0xF8FA: '薝' // U+859D <cjk>
	0xF8FB: '薟' // U+859F <cjk>
	0xF8FC: '𦿸' // U+26FF8 <cjk>
	0xF940: '𦿶' // U+26FF6 <cjk>
	0xF941: '𦿷' // U+26FF7 <cjk>
	0xF942: '薷' // U+85B7 <cjk>
	0xF943: '薼' // U+85BC <cjk>
	0xF944: '藇' // U+85C7 <cjk>
	0xF945: '藊' // U+85CA <cjk>
	0xF946: '藘' // U+85D8 <cjk>
	0xF947: '藙' // U+85D9 <cjk>
	0xF948: '藟' // U+85DF <cjk>
	0xF949: '藡' // U+85E1 <cjk>
	0xF94A: '藦' // U+85E6 <cjk>
	0xF94B: '藶' // U+85F6 <cjk>
	0xF94C: '蘀' // U+8600 <cjk>
	0xF94D: '蘑' // U+8611 <cjk>
	0xF94E: '蘞' // U+861E <cjk>
	0xF94F: '蘡' // U+8621 <cjk>
	0xF950: '蘤' // U+8624 <cjk>
	0xF951: '蘧' // U+8627 <cjk>
	0xF952: '𧄍' // U+2710D <cjk>
	0xF953: '蘹' // U+8639 <cjk>
	0xF954: '蘼' // U+863C <cjk>
	0xF955: '𧄹' // U+27139 <cjk>
	0xF956: '虀' // U+8640 <cjk>
	0xF957: '蘒' // U+FA20 CJK COMPATIBILITY IDEOGRAPH-FA20
	0xF958: '虓' // U+8653 <cjk>
	0xF959: '虖' // U+8656 <cjk>
	0xF95A: '虯' // U+866F <cjk>
	0xF95B: '虷' // U+8677 <cjk>
	0xF95C: '虺' // U+867A <cjk>
	0xF95D: '蚇' // U+8687 <cjk>
	0xF95E: '蚉' // U+8689 <cjk>
	0xF95F: '蚍' // U+868D <cjk>
	0xF960: '蚑' // U+8691 <cjk>
	0xF961: '蚜' // U+869C <cjk>
	0xF962: '蚝' // U+869D <cjk>
	0xF963: '蚨' // U+86A8 <cjk>
	0xF964: '﨡' // U+FA21 CJK COMPATIBILITY IDEOGRAPH-FA21
	0xF965: '蚱' // U+86B1 <cjk>
	0xF966: '蚳' // U+86B3 <cjk>
	0xF967: '蛁' // U+86C1 <cjk>
	0xF968: '蛃' // U+86C3 <cjk>
	0xF969: '蛑' // U+86D1 <cjk>
	0xF96A: '蛕' // U+86D5 <cjk>
	0xF96B: '蛗' // U+86D7 <cjk>
	0xF96C: '蛣' // U+86E3 <cjk>
	0xF96D: '蛦' // U+86E6 <cjk>
	0xF96E: '䖸' // U+45B8 <cjk>
	0xF96F: '蜅' // U+8705 <cjk>
	0xF970: '蜇' // U+8707 <cjk>
	0xF971: '蜎' // U+870E <cjk>
	0xF972: '蜐' // U+8710 <cjk>
	0xF973: '蜓' // U+8713 <cjk>
	0xF974: '蜙' // U+8719 <cjk>
	0xF975: '蜟' // U+871F <cjk>
	0xF976: '蜡' // U+8721 <cjk>
	0xF977: '蜣' // U+8723 <cjk>
	0xF978: '蜱' // U+8731 <cjk>
	0xF979: '蜺' // U+873A <cjk>
	0xF97A: '蜾' // U+873E <cjk>
	0xF97B: '蝀' // U+8740 <cjk>
	0xF97C: '蝃' // U+8743 <cjk>
	0xF97D: '蝑' // U+8751 <cjk>
	0xF97E: '蝘' // U+8758 <cjk>
	0xF980: '蝤' // U+8764 <cjk>
	0xF981: '蝥' // U+8765 <cjk>
	0xF982: '蝲' // U+8772 <cjk>
	0xF983: '蝼' // U+877C <cjk>
	0xF984: '𧏛' // U+273DB <cjk>
	0xF985: '𧏚' // U+273DA <cjk>
	0xF986: '螧' // U+87A7 <cjk>
	0xF987: '螉' // U+8789 <cjk>
	0xF988: '螋' // U+878B <cjk>
	0xF989: '螓' // U+8793 <cjk>
	0xF98A: '螠' // U+87A0 <cjk>
	0xF98B: '𧏾' // U+273FE <cjk>
	0xF98C: '䗥' // U+45E5 <cjk>
	0xF98D: '螾' // U+87BE <cjk>
	0xF98E: '𧐐' // U+27410 <cjk>
	0xF98F: '蟁' // U+87C1 <cjk>
	0xF990: '蟎' // U+87CE <cjk>
	0xF991: '蟵' // U+87F5 <cjk>
	0xF992: '蟟' // U+87DF <cjk>
	0xF993: '𧑉' // U+27449 <cjk>
	0xF994: '蟣' // U+87E3 <cjk>
	0xF995: '蟥' // U+87E5 <cjk>
	0xF996: '蟦' // U+87E6 <cjk>
	0xF997: '蟪' // U+87EA <cjk>
	0xF998: '蟫' // U+87EB <cjk>
	0xF999: '蟭' // U+87ED <cjk>
	0xF99A: '蠁' // U+8801 <cjk>
	0xF99B: '蠃' // U+8803 <cjk>
	0xF99C: '蠋' // U+880B <cjk>
	0xF99D: '蠓' // U+8813 <cjk>
	0xF99E: '蠨' // U+8828 <cjk>
	0xF99F: '蠮' // U+882E <cjk>
	0xF9A0: '蠲' // U+8832 <cjk>
	0xF9A1: '蠼' // U+883C <cjk>
	0xF9A2: '䘏' // U+460F <cjk>
	0xF9A3: '衊' // U+884A <cjk>
	0xF9A4: '衘' // U+8858 <cjk>
	0xF9A5: '衟' // U+885F <cjk>
	0xF9A6: '衤' // U+8864 <cjk>
	0xF9A7: '𧘕' // U+27615 <cjk>
	0xF9A8: '𧘔' // U+27614 <cjk>
	0xF9A9: '衩' // U+8869 <cjk>
	0xF9AA: '𧘱' // U+27631 <cjk>
	0xF9AB: '衯' // U+886F <cjk>
	0xF9AC: '袠' // U+88A0 <cjk>
	0xF9AD: '袼' // U+88BC <cjk>
	0xF9AE: '袽' // U+88BD <cjk>
	0xF9AF: '袾' // U+88BE <cjk>
	0xF9B0: '裀' // U+88C0 <cjk>
	0xF9B1: '裒' // U+88D2 <cjk>
	0xF9B2: '𧚓' // U+27693 <cjk>
	0xF9B3: '裑' // U+88D1 <cjk>
	0xF9B4: '裓' // U+88D3 <cjk>
	0xF9B5: '裛' // U+88DB <cjk>
	0xF9B6: '裰' // U+88F0 <cjk>
	0xF9B7: '裱' // U+88F1 <cjk>
	0xF9B8: '䙁' // U+4641 <cjk>
	0xF9B9: '褁' // U+8901 <cjk>
	0xF9BA: '𧜎' // U+2770E <cjk>
	0xF9BB: '褷' // U+8937 <cjk>
	0xF9BC: '𧜣' // U+27723 <cjk>
	0xF9BD: '襂' // U+8942 <cjk>
	0xF9BE: '襅' // U+8945 <cjk>
	0xF9BF: '襉' // U+8949 <cjk>
	0xF9C0: '𧝒' // U+27752 <cjk>
	0xF9C1: '䙥' // U+4665 <cjk>
	0xF9C2: '襢' // U+8962 <cjk>
	0xF9C3: '覀' // U+8980 <cjk>
	0xF9C4: '覉' // U+8989 <cjk>
	0xF9C5: '覐' // U+8990 <cjk>
	0xF9C6: '覟' // U+899F <cjk>
	0xF9C7: '覰' // U+89B0 <cjk>
	0xF9C8: '覷' // U+89B7 <cjk>
	0xF9C9: '觖' // U+89D6 <cjk>
	0xF9CA: '觘' // U+89D8 <cjk>
	0xF9CB: '觫' // U+89EB <cjk>
	0xF9CC: '䚡' // U+46A1 <cjk>
	0xF9CD: '觱' // U+89F1 <cjk>
	0xF9CE: '觳' // U+89F3 <cjk>
	0xF9CF: '觽' // U+89FD <cjk>
	0xF9D0: '觿' // U+89FF <cjk>
	0xF9D1: '䚯' // U+46AF <cjk>
	0xF9D2: '訑' // U+8A11 <cjk>
	0xF9D3: '訔' // U+8A14 <cjk>
	0xF9D4: '𧦅' // U+27985 <cjk>
	0xF9D5: '訡' // U+8A21 <cjk>
	0xF9D6: '訵' // U+8A35 <cjk>
	0xF9D7: '訾' // U+8A3E <cjk>
	0xF9D8: '詅' // U+8A45 <cjk>
	0xF9D9: '詍' // U+8A4D <cjk>
	0xF9DA: '詘' // U+8A58 <cjk>
	0xF9DB: '誮' // U+8AAE <cjk>
	0xF9DC: '誐' // U+8A90 <cjk>
	0xF9DD: '誷' // U+8AB7 <cjk>
	0xF9DE: '誾' // U+8ABE <cjk>
	0xF9DF: '諗' // U+8AD7 <cjk>
	0xF9E0: '諼' // U+8AFC <cjk>
	0xF9E1: '𧪄' // U+27A84 <cjk>
	0xF9E2: '謊' // U+8B0A <cjk>
	0xF9E3: '謅' // U+8B05 <cjk>
	0xF9E4: '謍' // U+8B0D <cjk>
	0xF9E5: '謜' // U+8B1C <cjk>
	0xF9E6: '謟' // U+8B1F <cjk>
	0xF9E7: '謭' // U+8B2D <cjk>
	0xF9E8: '譃' // U+8B43 <cjk>
	0xF9E9: '䜌' // U+470C <cjk>
	0xF9EA: '譑' // U+8B51 <cjk>
	0xF9EB: '譞' // U+8B5E <cjk>
	0xF9EC: '譶' // U+8B76 <cjk>
	0xF9ED: '譿' // U+8B7F <cjk>
	0xF9EE: '讁' // U+8B81 <cjk>
	0xF9EF: '讋' // U+8B8B <cjk>
	0xF9F0: '讔' // U+8B94 <cjk>
	0xF9F1: '讕' // U+8B95 <cjk>
	0xF9F2: '讜' // U+8B9C <cjk>
	0xF9F3: '讞' // U+8B9E <cjk>
	0xF9F4: '谹' // U+8C39 <cjk>
	0xF9F5: '𧮳' // U+27BB3 <cjk>
	0xF9F6: '谽' // U+8C3D <cjk>
	0xF9F7: '𧮾' // U+27BBE <cjk>
	0xF9F8: '𧯇' // U+27BC7 <cjk>
	0xF9F9: '豅' // U+8C45 <cjk>
	0xF9FA: '豇' // U+8C47 <cjk>
	0xF9FB: '豏' // U+8C4F <cjk>
	0xF9FC: '豔' // U+8C54 <cjk>
	0xFA40: '豗' // U+8C57 <cjk>
	0xFA41: '豩' // U+8C69 <cjk>
	0xFA42: '豭' // U+8C6D <cjk>
	0xFA43: '豳' // U+8C73 <cjk>
	0xFA44: '𧲸' // U+27CB8 <cjk>
	0xFA45: '貓' // U+8C93 <cjk>
	0xFA46: '貒' // U+8C92 <cjk>
	0xFA47: '貙' // U+8C99 <cjk>
	0xFA48: '䝤' // U+4764 <cjk>
	0xFA49: '貛' // U+8C9B <cjk>
	0xFA4A: '貤' // U+8CA4 <cjk>
	0xFA4B: '賖' // U+8CD6 <cjk>
	0xFA4C: '賕' // U+8CD5 <cjk>
	0xFA4D: '賙' // U+8CD9 <cjk>
	0xFA4E: '𧶠' // U+27DA0 <cjk>
	0xFA4F: '賰' // U+8CF0 <cjk>
	0xFA50: '賱' // U+8CF1 <cjk>
	0xFA51: '𧸐' // U+27E10 <cjk>
	0xFA52: '贉' // U+8D09 <cjk>
	0xFA53: '贎' // U+8D0E <cjk>
	0xFA54: '赬' // U+8D6C <cjk>
	0xFA55: '趄' // U+8D84 <cjk>
	0xFA56: '趕' // U+8D95 <cjk>
	0xFA57: '趦' // U+8DA6 <cjk>
	0xFA58: '𧾷' // U+27FB7 <cjk>
	0xFA59: '跆' // U+8DC6 <cjk>
	0xFA5A: '跈' // U+8DC8 <cjk>
	0xFA5B: '跙' // U+8DD9 <cjk>
	0xFA5C: '跬' // U+8DEC <cjk>
	0xFA5D: '踌' // U+8E0C <cjk>
	0xFA5E: '䟽' // U+47FD <cjk>
	0xFA5F: '跽' // U+8DFD <cjk>
	0xFA60: '踆' // U+8E06 <cjk>
	0xFA61: '𨂊' // U+2808A <cjk>
	0xFA62: '踔' // U+8E14 <cjk>
	0xFA63: '踖' // U+8E16 <cjk>
	0xFA64: '踡' // U+8E21 <cjk>
	0xFA65: '踢' // U+8E22 <cjk>
	0xFA66: '踧' // U+8E27 <cjk>
	0xFA67: '𨂻' // U+280BB <cjk>
	0xFA68: '䠖' // U+4816 <cjk>
	0xFA69: '踶' // U+8E36 <cjk>
	0xFA6A: '踹' // U+8E39 <cjk>
	0xFA6B: '蹋' // U+8E4B <cjk>
	0xFA6C: '蹔' // U+8E54 <cjk>
	0xFA6D: '蹢' // U+8E62 <cjk>
	0xFA6E: '蹬' // U+8E6C <cjk>
	0xFA6F: '蹭' // U+8E6D <cjk>
	0xFA70: '蹯' // U+8E6F <cjk>
	0xFA71: '躘' // U+8E98 <cjk>
	0xFA72: '躞' // U+8E9E <cjk>
	0xFA73: '躮' // U+8EAE <cjk>
	0xFA74: '躳' // U+8EB3 <cjk>
	0xFA75: '躵' // U+8EB5 <cjk>
	0xFA76: '躶' // U+8EB6 <cjk>
	0xFA77: '躻' // U+8EBB <cjk>
	0xFA78: '𨊂' // U+28282 <cjk>
	0xFA79: '軑' // U+8ED1 <cjk>
	0xFA7A: '軔' // U+8ED4 <cjk>
	0xFA7B: '䡎' // U+484E <cjk>
	0xFA7C: '軹' // U+8EF9 <cjk>
	0xFA7D: '𨋳' // U+282F3 <cjk>
	0xFA7E: '輀' // U+8F00 <cjk>
	0xFA80: '輈' // U+8F08 <cjk>
	0xFA81: '輗' // U+8F17 <cjk>
	0xFA82: '輫' // U+8F2B <cjk>
	0xFA83: '轀' // U+8F40 <cjk>
	0xFA84: '轊' // U+8F4A <cjk>
	0xFA85: '轘' // U+8F58 <cjk>
	0xFA86: '𨐌' // U+2840C <cjk>
	0xFA87: '辤' // U+8FA4 <cjk>
	0xFA88: '辴' // U+8FB4 <cjk>
	0xFA89: '辶' // U+FA66 CJK COMPATIBILITY IDEOGRAPH-FA66
	0xFA8A: '辶' // U+8FB6 <cjk>
	0xFA8B: '𨑕' // U+28455 <cjk>
	0xFA8C: '迁' // U+8FC1 <cjk>
	0xFA8D: '迆' // U+8FC6 <cjk>
	0xFA8E: '﨤' // U+FA24 CJK COMPATIBILITY IDEOGRAPH-FA24
	0xFA8F: '迊' // U+8FCA <cjk>
	0xFA90: '迍' // U+8FCD <cjk>
	0xFA91: '迓' // U+8FD3 <cjk>
	0xFA92: '迕' // U+8FD5 <cjk>
	0xFA93: '迠' // U+8FE0 <cjk>
	0xFA94: '迱' // U+8FF1 <cjk>
	0xFA95: '迵' // U+8FF5 <cjk>
	0xFA96: '迻' // U+8FFB <cjk>
	0xFA97: '适' // U+9002 <cjk>
	0xFA98: '逌' // U+900C <cjk>
	0xFA99: '逷' // U+9037 <cjk>
	0xFA9A: '𨕫' // U+2856B <cjk>
	0xFA9B: '遃' // U+9043 <cjk>
	0xFA9C: '遄' // U+9044 <cjk>
	0xFA9D: '遝' // U+905D <cjk>
	0xFA9E: '𨗈' // U+285C8 <cjk>
	0xFA9F: '𨗉' // U+285C9 <cjk>
	0xFAA0: '邅' // U+9085 <cjk>
	0xFAA1: '邌' // U+908C <cjk>
	0xFAA2: '邐' // U+9090 <cjk>
	0xFAA3: '阝' // U+961D <cjk>
	0xFAA4: '邡' // U+90A1 <cjk>
	0xFAA5: '䢵' // U+48B5 <cjk>
	0xFAA6: '邰' // U+90B0 <cjk>
	0xFAA7: '邶' // U+90B6 <cjk>
	0xFAA8: '郃' // U+90C3 <cjk>
	0xFAA9: '郈' // U+90C8 <cjk>
	0xFAAA: '𨛗' // U+286D7 <cjk>
	0xFAAB: '郜' // U+90DC <cjk>
	0xFAAC: '郟' // U+90DF <cjk>
	0xFAAD: '𨛺' // U+286FA <cjk>
	0xFAAE: '郶' // U+90F6 <cjk>
	0xFAAF: '郲' // U+90F2 <cjk>
	0xFAB0: '鄀' // U+9100 <cjk>
	0xFAB1: '郫' // U+90EB <cjk>
	0xFAB2: '郾' // U+90FE <cjk>
	0xFAB3: '郿' // U+90FF <cjk>
	0xFAB4: '鄄' // U+9104 <cjk>
	0xFAB5: '鄆' // U+9106 <cjk>
	0xFAB6: '鄘' // U+9118 <cjk>
	0xFAB7: '鄜' // U+911C <cjk>
	0xFAB8: '鄞' // U+911E <cjk>
	0xFAB9: '鄷' // U+9137 <cjk>
	0xFABA: '鄹' // U+9139 <cjk>
	0xFABB: '鄺' // U+913A <cjk>
	0xFABC: '酆' // U+9146 <cjk>
	0xFABD: '酇' // U+9147 <cjk>
	0xFABE: '酗' // U+9157 <cjk>
	0xFABF: '酙' // U+9159 <cjk>
	0xFAC0: '酡' // U+9161 <cjk>
	0xFAC1: '酤' // U+9164 <cjk>
	0xFAC2: '酴' // U+9174 <cjk>
	0xFAC3: '酹' // U+9179 <cjk>
	0xFAC4: '醅' // U+9185 <cjk>
	0xFAC5: '醎' // U+918E <cjk>
	0xFAC6: '醨' // U+91A8 <cjk>
	0xFAC7: '醮' // U+91AE <cjk>
	0xFAC8: '醳' // U+91B3 <cjk>
	0xFAC9: '醶' // U+91B6 <cjk>
	0xFACA: '釃' // U+91C3 <cjk>
	0xFACB: '釄' // U+91C4 <cjk>
	0xFACC: '釚' // U+91DA <cjk>
	0xFACD: '𨥉' // U+28949 <cjk>
	0xFACE: '𨥆' // U+28946 <cjk>
	0xFACF: '釬' // U+91EC <cjk>
	0xFAD0: '釮' // U+91EE <cjk>
	0xFAD1: '鈁' // U+9201 <cjk>
	0xFAD2: '鈊' // U+920A <cjk>
	0xFAD3: '鈖' // U+9216 <cjk>
	0xFAD4: '鈗' // U+9217 <cjk>
	0xFAD5: '𨥫' // U+2896B <cjk>
	0xFAD6: '鈳' // U+9233 <cjk>
	0xFAD7: '鉂' // U+9242 <cjk>
	0xFAD8: '鉇' // U+9247 <cjk>
	0xFAD9: '鉊' // U+924A <cjk>
	0xFADA: '鉎' // U+924E <cjk>
	0xFADB: '鉑' // U+9251 <cjk>
	0xFADC: '鉖' // U+9256 <cjk>
	0xFADD: '鉙' // U+9259 <cjk>
	0xFADE: '鉠' // U+9260 <cjk>
	0xFADF: '鉡' // U+9261 <cjk>
	0xFAE0: '鉥' // U+9265 <cjk>
	0xFAE1: '鉧' // U+9267 <cjk>
	0xFAE2: '鉨' // U+9268 <cjk>
	0xFAE3: '𨦇' // U+28987 <cjk>
	0xFAE4: '𨦈' // U+28988 <cjk>
	0xFAE5: '鉼' // U+927C <cjk>
	0xFAE6: '鉽' // U+927D <cjk>
	0xFAE7: '鉿' // U+927F <cjk>
	0xFAE8: '銉' // U+9289 <cjk>
	0xFAE9: '銍' // U+928D <cjk>
	0xFAEA: '銗' // U+9297 <cjk>
	0xFAEB: '銙' // U+9299 <cjk>
	0xFAEC: '銟' // U+929F <cjk>
	0xFAED: '銧' // U+92A7 <cjk>
	0xFAEE: '銫' // U+92AB <cjk>
	0xFAEF: '𨦺' // U+289BA <cjk>
	0xFAF0: '𨦻' // U+289BB <cjk>
	0xFAF1: '銲' // U+92B2 <cjk>
	0xFAF2: '銿' // U+92BF <cjk>
	0xFAF3: '鋀' // U+92C0 <cjk>
	0xFAF4: '鋆' // U+92C6 <cjk>
	0xFAF5: '鋎' // U+92CE <cjk>
	0xFAF6: '鋐' // U+92D0 <cjk>
	0xFAF7: '鋗' // U+92D7 <cjk>
	0xFAF8: '鋙' // U+92D9 <cjk>
	0xFAF9: '鋥' // U+92E5 <cjk>
	0xFAFA: '鋧' // U+92E7 <cjk>
	0xFAFB: '錑' // U+9311 <cjk>
	0xFAFC: '𨨞' // U+28A1E <cjk>
	0xFB40: '𨨩' // U+28A29 <cjk>
	0xFB41: '鋷' // U+92F7 <cjk>
	0xFB42: '鋹' // U+92F9 <cjk>
	0xFB43: '鋻' // U+92FB <cjk>
	0xFB44: '錂' // U+9302 <cjk>
	0xFB45: '錍' // U+930D <cjk>
	0xFB46: '錕' // U+9315 <cjk>
	0xFB47: '錝' // U+931D <cjk>
	0xFB48: '錞' // U+931E <cjk>
	0xFB49: '錧' // U+9327 <cjk>
	0xFB4A: '錩' // U+9329 <cjk>
	0xFB4B: '𨩱' // U+28A71 <cjk>
	0xFB4C: '𨩃' // U+28A43 <cjk>
	0xFB4D: '鍇' // U+9347 <cjk>
	0xFB4E: '鍑' // U+9351 <cjk>
	0xFB4F: '鍗' // U+9357 <cjk>
	0xFB50: '鍚' // U+935A <cjk>
	0xFB51: '鍫' // U+936B <cjk>
	0xFB52: '鍱' // U+9371 <cjk>
	0xFB53: '鍳' // U+9373 <cjk>
	0xFB54: '鎡' // U+93A1 <cjk>
	0xFB55: '𨪙' // U+28A99 <cjk>
	0xFB56: '𨫍' // U+28ACD <cjk>
	0xFB57: '鎈' // U+9388 <cjk>
	0xFB58: '鎋' // U+938B <cjk>
	0xFB59: '鎏' // U+938F <cjk>
	0xFB5A: '鎞' // U+939E <cjk>
	0xFB5B: '鏵' // U+93F5 <cjk>
	0xFB5C: '𨫤' // U+28AE4 <cjk>
	0xFB5D: '𨫝' // U+28ADD <cjk>
	0xFB5E: '鏱' // U+93F1 <cjk>
	0xFB5F: '鏁' // U+93C1 <cjk>
	0xFB60: '鏇' // U+93C7 <cjk>
	0xFB61: '鏜' // U+93DC <cjk>
	0xFB62: '鏢' // U+93E2 <cjk>
	0xFB63: '鏧' // U+93E7 <cjk>
	0xFB64: '鐉' // U+9409 <cjk>
	0xFB65: '鐏' // U+940F <cjk>
	0xFB66: '鐖' // U+9416 <cjk>
	0xFB67: '鐗' // U+9417 <cjk>
	0xFB68: '鏻' // U+93FB <cjk>
	0xFB69: '鐲' // U+9432 <cjk>
	0xFB6A: '鐴' // U+9434 <cjk>
	0xFB6B: '鐻' // U+943B <cjk>
	0xFB6C: '鑅' // U+9445 <cjk>
	0xFB6D: '𨯁' // U+28BC1 <cjk>
	0xFB6E: '𨯯' // U+28BEF <cjk>
	0xFB6F: '鑭' // U+946D <cjk>
	0xFB70: '鑯' // U+946F <cjk>
	0xFB71: '镸' // U+9578 <cjk>
	0xFB72: '镹' // U+9579 <cjk>
	0xFB73: '閆' // U+9586 <cjk>
	0xFB74: '閌' // U+958C <cjk>
	0xFB75: '閍' // U+958D <cjk>
	0xFB76: '𨴐' // U+28D10 <cjk>
	0xFB77: '閫' // U+95AB <cjk>
	0xFB78: '閴' // U+95B4 <cjk>
	0xFB79: '𨵱' // U+28D71 <cjk>
	0xFB7A: '闈' // U+95C8 <cjk>
	0xFB7B: '𨷻' // U+28DFB <cjk>
	0xFB7C: '𨸟' // U+28E1F <cjk>
	0xFB7D: '阬' // U+962C <cjk>
	0xFB7E: '阳' // U+9633 <cjk>
	0xFB80: '阴' // U+9634 <cjk>
	0xFB81: '𨸶' // U+28E36 <cjk>
	0xFB82: '阼' // U+963C <cjk>
	0xFB83: '陁' // U+9641 <cjk>
	0xFB84: '陡' // U+9661 <cjk>
	0xFB85: '𨺉' // U+28E89 <cjk>
	0xFB86: '隂' // U+9682 <cjk>
	0xFB87: '𨻫' // U+28EEB <cjk>
	0xFB88: '隚' // U+969A <cjk>
	0xFB89: '𨼲' // U+28F32 <cjk>
	0xFB8A: '䧧' // U+49E7 <cjk>
	0xFB8B: '隩' // U+96A9 <cjk>
	0xFB8C: '隯' // U+96AF <cjk>
	0xFB8D: '隳' // U+96B3 <cjk>
	0xFB8E: '隺' // U+96BA <cjk>
	0xFB8F: '隽' // U+96BD <cjk>
	0xFB90: '䧺' // U+49FA <cjk>
	0xFB91: '𨿸' // U+28FF8 <cjk>
	0xFB92: '雘' // U+96D8 <cjk>
	0xFB93: '雚' // U+96DA <cjk>
	0xFB94: '雝' // U+96DD <cjk>
	0xFB95: '䨄' // U+4A04 <cjk>
	0xFB96: '霔' // U+9714 <cjk>
	0xFB97: '霣' // U+9723 <cjk>
	0xFB98: '䨩' // U+4A29 <cjk>
	0xFB99: '霶' // U+9736 <cjk>
	0xFB9A: '靁' // U+9741 <cjk>
	0xFB9B: '靇' // U+9747 <cjk>
	0xFB9C: '靕' // U+9755 <cjk>
	0xFB9D: '靗' // U+9757 <cjk>
	0xFB9E: '靛' // U+975B <cjk>
	0xFB9F: '靪' // U+976A <cjk>
	0xFBA0: '𩊠' // U+292A0 <cjk>
	0xFBA1: '𩊱' // U+292B1 <cjk>
	0xFBA2: '鞖' // U+9796 <cjk>
	0xFBA3: '鞚' // U+979A <cjk>
	0xFBA4: '鞞' // U+979E <cjk>
	0xFBA5: '鞢' // U+97A2 <cjk>
	0xFBA6: '鞱' // U+97B1 <cjk>
	0xFBA7: '鞲' // U+97B2 <cjk>
	0xFBA8: '鞾' // U+97BE <cjk>
	0xFBA9: '韌' // U+97CC <cjk>
	0xFBAA: '韑' // U+97D1 <cjk>
	0xFBAB: '韔' // U+97D4 <cjk>
	0xFBAC: '韘' // U+97D8 <cjk>
	0xFBAD: '韙' // U+97D9 <cjk>
	0xFBAE: '韡' // U+97E1 <cjk>
	0xFBAF: '韱' // U+97F1 <cjk>
	0xFBB0: '頄' // U+9804 <cjk>
	0xFBB1: '頍' // U+980D <cjk>
	0xFBB2: '頎' // U+980E <cjk>
	0xFBB3: '頔' // U+9814 <cjk>
	0xFBB4: '頖' // U+9816 <cjk>
	0xFBB5: '䪼' // U+4ABC <cjk>
	0xFBB6: '𩒐' // U+29490 <cjk>
	0xFBB7: '頣' // U+9823 <cjk>
	0xFBB8: '頲' // U+9832 <cjk>
	0xFBB9: '頳' // U+9833 <cjk>
	0xFBBA: '頥' // U+9825 <cjk>
	0xFBBB: '顇' // U+9847 <cjk>
	0xFBBC: '顦' // U+9866 <cjk>
	0xFBBD: '颫' // U+98AB <cjk>
	0xFBBE: '颭' // U+98AD <cjk>
	0xFBBF: '颰' // U+98B0 <cjk>
	0xFBC0: '𩗏' // U+295CF <cjk>
	0xFBC1: '颷' // U+98B7 <cjk>
	0xFBC2: '颸' // U+98B8 <cjk>
	0xFBC3: '颻' // U+98BB <cjk>
	0xFBC4: '颼' // U+98BC <cjk>
	0xFBC5: '颿' // U+98BF <cjk>
	0xFBC6: '飂' // U+98C2 <cjk>
	0xFBC7: '飇' // U+98C7 <cjk>
	0xFBC8: '飋' // U+98CB <cjk>
	0xFBC9: '飠' // U+98E0 <cjk>
	0xFBCA: '𩙿' // U+2967F <cjk>
	0xFBCB: '飡' // U+98E1 <cjk>
	0xFBCC: '飣' // U+98E3 <cjk>
	0xFBCD: '飥' // U+98E5 <cjk>
	0xFBCE: '飪' // U+98EA <cjk>
	0xFBCF: '飰' // U+98F0 <cjk>
	0xFBD0: '飱' // U+98F1 <cjk>
	0xFBD1: '飳' // U+98F3 <cjk>
	0xFBD2: '餈' // U+9908 <cjk>
	0xFBD3: '䬻' // U+4B3B <cjk>
	0xFBD4: '𩛰' // U+296F0 <cjk>
	0xFBD5: '餖' // U+9916 <cjk>
	0xFBD6: '餗' // U+9917 <cjk>
	0xFBD7: '𩜙' // U+29719 <cjk>
	0xFBD8: '餚' // U+991A <cjk>
	0xFBD9: '餛' // U+991B <cjk>
	0xFBDA: '餜' // U+991C <cjk>
	0xFBDB: '𩝐' // U+29750 <cjk>
	0xFBDC: '餱' // U+9931 <cjk>
	0xFBDD: '餲' // U+9932 <cjk>
	0xFBDE: '餳' // U+9933 <cjk>
	0xFBDF: '餺' // U+993A <cjk>
	0xFBE0: '餻' // U+993B <cjk>
	0xFBE1: '餼' // U+993C <cjk>
	0xFBE2: '饀' // U+9940 <cjk>
	0xFBE3: '饁' // U+9941 <cjk>
	0xFBE4: '饆' // U+9946 <cjk>
	0xFBE5: '饍' // U+994D <cjk>
	0xFBE6: '饎' // U+994E <cjk>
	0xFBE7: '饜' // U+995C <cjk>
	0xFBE8: '饟' // U+995F <cjk>
	0xFBE9: '饠' // U+9960 <cjk>
	0xFBEA: '馣' // U+99A3 <cjk>
	0xFBEB: '馦' // U+99A6 <cjk>
	0xFBEC: '馹' // U+99B9 <cjk>
	0xFBED: '馽' // U+99BD <cjk>
	0xFBEE: '馿' // U+99BF <cjk>
	0xFBEF: '駃' // U+99C3 <cjk>
	0xFBF0: '駉' // U+99C9 <cjk>
	0xFBF1: '駔' // U+99D4 <cjk>
	0xFBF2: '駙' // U+99D9 <cjk>
	0xFBF3: '駞' // U+99DE <cjk>
	0xFBF4: '𩣆' // U+298C6 <cjk>
	0xFBF5: '駰' // U+99F0 <cjk>
	0xFBF6: '駹' // U+99F9 <cjk>
	0xFBF7: '駼' // U+99FC <cjk>
	0xFBF8: '騊' // U+9A0A <cjk>
	0xFBF9: '騑' // U+9A11 <cjk>
	0xFBFA: '騖' // U+9A16 <cjk>
	0xFBFB: '騚' // U+9A1A <cjk>
	0xFBFC: '騠' // U+9A20 <cjk>
	0xFC40: '騱' // U+9A31 <cjk>
	0xFC41: '騶' // U+9A36 <cjk>
	0xFC42: '驄' // U+9A44 <cjk>
	0xFC43: '驌' // U+9A4C <cjk>
	0xFC44: '驘' // U+9A58 <cjk>
	0xFC45: '䯂' // U+4BC2 <cjk>
	0xFC46: '骯' // U+9AAF <cjk>
	0xFC47: '䯊' // U+4BCA <cjk>
	0xFC48: '骷' // U+9AB7 <cjk>
	0xFC49: '䯒' // U+4BD2 <cjk>
	0xFC4A: '骹' // U+9AB9 <cjk>
	0xFC4B: '𩩲' // U+29A72 <cjk>
	0xFC4C: '髆' // U+9AC6 <cjk>
	0xFC4D: '髐' // U+9AD0 <cjk>
	0xFC4E: '髒' // U+9AD2 <cjk>
	0xFC4F: '髕' // U+9AD5 <cjk>
	0xFC50: '䯨' // U+4BE8 <cjk>
	0xFC51: '髜' // U+9ADC <cjk>
	0xFC52: '髠' // U+9AE0 <cjk>
	0xFC53: '髥' // U+9AE5 <cjk>
	0xFC54: '髩' // U+9AE9 <cjk>
	0xFC55: '鬃' // U+9B03 <cjk>
	0xFC56: '鬌' // U+9B0C <cjk>
	0xFC57: '鬐' // U+9B10 <cjk>
	0xFC58: '鬒' // U+9B12 <cjk>
	0xFC59: '鬖' // U+9B16 <cjk>
	0xFC5A: '鬜' // U+9B1C <cjk>
	0xFC5B: '鬫' // U+9B2B <cjk>
	0xFC5C: '鬳' // U+9B33 <cjk>
	0xFC5D: '鬽' // U+9B3D <cjk>
	0xFC5E: '䰠' // U+4C20 <cjk>
	0xFC5F: '魋' // U+9B4B <cjk>
	0xFC60: '魣' // U+9B63 <cjk>
	0xFC61: '魥' // U+9B65 <cjk>
	0xFC62: '魫' // U+9B6B <cjk>
	0xFC63: '魬' // U+9B6C <cjk>
	0xFC64: '魳' // U+9B73 <cjk>
	0xFC65: '魶' // U+9B76 <cjk>
	0xFC66: '魷' // U+9B77 <cjk>
	0xFC67: '鮦' // U+9BA6 <cjk>
	0xFC68: '鮬' // U+9BAC <cjk>
	0xFC69: '鮱' // U+9BB1 <cjk>
	0xFC6A: '𩷛' // U+29DDB <cjk>
	0xFC6B: '𩸽' // U+29E3D <cjk>
	0xFC6C: '鮲' // U+9BB2 <cjk>
	0xFC6D: '鮸' // U+9BB8 <cjk>
	0xFC6E: '鮾' // U+9BBE <cjk>
	0xFC6F: '鯇' // U+9BC7 <cjk>
	0xFC70: '鯳' // U+9BF3 <cjk>
	0xFC71: '鯘' // U+9BD8 <cjk>
	0xFC72: '鯝' // U+9BDD <cjk>
	0xFC73: '鯧' // U+9BE7 <cjk>
	0xFC74: '鯪' // U+9BEA <cjk>
	0xFC75: '鯫' // U+9BEB <cjk>
	0xFC76: '鯯' // U+9BEF <cjk>
	0xFC77: '鯮' // U+9BEE <cjk>
	0xFC78: '𩸕' // U+29E15 <cjk>
	0xFC79: '鯺' // U+9BFA <cjk>
	0xFC7A: '𩺊' // U+29E8A <cjk>
	0xFC7B: '鯷' // U+9BF7 <cjk>
	0xFC7C: '𩹉' // U+29E49 <cjk>
	0xFC7D: '鰖' // U+9C16 <cjk>
	0xFC7E: '鰘' // U+9C18 <cjk>
	0xFC80: '鰙' // U+9C19 <cjk>
	0xFC81: '鰚' // U+9C1A <cjk>
	0xFC82: '鰝' // U+9C1D <cjk>
	0xFC83: '鰢' // U+9C22 <cjk>
	0xFC84: '鰧' // U+9C27 <cjk>
	0xFC85: '鰩' // U+9C29 <cjk>
	0xFC86: '鰪' // U+9C2A <cjk>
	0xFC87: '𩻄' // U+29EC4 <cjk>
	0xFC88: '鰱' // U+9C31 <cjk>
	0xFC89: '鰶' // U+9C36 <cjk>
	0xFC8A: '鰷' // U+9C37 <cjk>
	0xFC8B: '鱅' // U+9C45 <cjk>
	0xFC8C: '鱜' // U+9C5C <cjk>
	0xFC8D: '𩻩' // U+29EE9 <cjk>
	0xFC8E: '鱉' // U+9C49 <cjk>
	0xFC8F: '鱊' // U+9C4A <cjk>
	0xFC90: '𩻛' // U+29EDB <cjk>
	0xFC91: '鱔' // U+9C54 <cjk>
	0xFC92: '鱘' // U+9C58 <cjk>
	0xFC93: '鱛' // U+9C5B <cjk>
	0xFC94: '鱝' // U+9C5D <cjk>
	0xFC95: '鱟' // U+9C5F <cjk>
	0xFC96: '鱩' // U+9C69 <cjk>
	0xFC97: '鱪' // U+9C6A <cjk>
	0xFC98: '鱫' // U+9C6B <cjk>
	0xFC99: '鱭' // U+9C6D <cjk>
	0xFC9A: '鱮' // U+9C6E <cjk>
	0xFC9B: '鱰' // U+9C70 <cjk>
	0xFC9C: '鱲' // U+9C72 <cjk>
	0xFC9D: '鱵' // U+9C75 <cjk>
	0xFC9E: '鱺' // U+9C7A <cjk>
	0xFC9F: '鳦' // U+9CE6 <cjk>
	0xFCA0: '鳲' // U+9CF2 <cjk>
	0xFCA1: '鴋' // U+9D0B <cjk>
	0xFCA2: '鴂' // U+9D02 <cjk>
	0xFCA3: '𩿎' // U+29FCE <cjk>
	0xFCA4: '鴑' // U+9D11 <cjk>
	0xFCA5: '鴗' // U+9D17 <cjk>
	0xFCA6: '鴘' // U+9D18 <cjk>
	0xFCA7: '𪀯' // U+2A02F <cjk>
	0xFCA8: '䳄' // U+4CC4 <cjk>
	0xFCA9: '𪀚' // U+2A01A <cjk>
	0xFCAA: '鴲' // U+9D32 <cjk>
	0xFCAB: '䳑' // U+4CD1 <cjk>
	0xFCAC: '鵂' // U+9D42 <cjk>
	0xFCAD: '鵊' // U+9D4A <cjk>
	0xFCAE: '鵟' // U+9D5F <cjk>
	0xFCAF: '鵢' // U+9D62 <cjk>
	0xFCB0: '𪃹' // U+2A0F9 <cjk>
	0xFCB1: '鵩' // U+9D69 <cjk>
	0xFCB2: '鵫' // U+9D6B <cjk>
	0xFCB3: '𪂂' // U+2A082 <cjk>
	0xFCB4: '鵳' // U+9D73 <cjk>
	0xFCB5: '鵶' // U+9D76 <cjk>
	0xFCB6: '鵷' // U+9D77 <cjk>
	0xFCB7: '鵾' // U+9D7E <cjk>
	0xFCB8: '鶄' // U+9D84 <cjk>
	0xFCB9: '鶍' // U+9D8D <cjk>
	0xFCBA: '鶙' // U+9D99 <cjk>
	0xFCBB: '鶡' // U+9DA1 <cjk>
	0xFCBC: '鶿' // U+9DBF <cjk>
	0xFCBD: '鶵' // U+9DB5 <cjk>
	0xFCBE: '鶹' // U+9DB9 <cjk>
	0xFCBF: '鶽' // U+9DBD <cjk>
	0xFCC0: '鷃' // U+9DC3 <cjk>
	0xFCC1: '鷇' // U+9DC7 <cjk>
	0xFCC2: '鷉' // U+9DC9 <cjk>
	0xFCC3: '鷖' // U+9DD6 <cjk>
	0xFCC4: '鷚' // U+9DDA <cjk>
	0xFCC5: '鷟' // U+9DDF <cjk>
	0xFCC6: '鷠' // U+9DE0 <cjk>
	0xFCC7: '鷣' // U+9DE3 <cjk>
	0xFCC8: '鷴' // U+9DF4 <cjk>
	0xFCC9: '䴇' // U+4D07 <cjk>
	0xFCCA: '鸊' // U+9E0A <cjk>
	0xFCCB: '鸂' // U+9E02 <cjk>
	0xFCCC: '鸍' // U+9E0D <cjk>
	0xFCCD: '鸙' // U+9E19 <cjk>
	0xFCCE: '鸜' // U+9E1C <cjk>
	0xFCCF: '鸝' // U+9E1D <cjk>
	0xFCD0: '鹻' // U+9E7B <cjk>
	0xFCD1: '𢈘' // U+22218 <cjk>
	0xFCD2: '麀' // U+9E80 <cjk>
	0xFCD3: '麅' // U+9E85 <cjk>
	0xFCD4: '麛' // U+9E9B <cjk>
	0xFCD5: '麨' // U+9EA8 <cjk>
	0xFCD6: '𪎌' // U+2A38C <cjk>
	0xFCD7: '麽' // U+9EBD <cjk>
	0xFCD8: '𪐷' // U+2A437 <cjk>
	0xFCD9: '黟' // U+9EDF <cjk>
	0xFCDA: '黧' // U+9EE7 <cjk>
	0xFCDB: '黮' // U+9EEE <cjk>
	0xFCDC: '黿' // U+9EFF <cjk>
	0xFCDD: '鼂' // U+9F02 <cjk>
	0xFCDE: '䵷' // U+4D77 <cjk>
	0xFCDF: '鼃' // U+9F03 <cjk>
	0xFCE0: '鼗' // U+9F17 <cjk>
	0xFCE1: '鼙' // U+9F19 <cjk>
	0xFCE2: '鼯' // U+9F2F <cjk>
	0xFCE3: '鼷' // U+9F37 <cjk>
	0xFCE4: '鼺' // U+9F3A <cjk>
	0xFCE5: '鼽' // U+9F3D <cjk>
	0xFCE6: '齁' // U+9F41 <cjk>
	0xFCE7: '齅' // U+9F45 <cjk>
	0xFCE8: '齆' // U+9F46 <cjk>
	0xFCE9: '齓' // U+9F53 <cjk>
	0xFCEA: '齕' // U+9F55 <cjk>
	0xFCEB: '齘' // U+9F58 <cjk>
	0xFCEC: '𪗱' // U+2A5F1 <cjk>
	0xFCED: '齝' // U+9F5D <cjk>
	0xFCEE: '𪘂' // U+2A602 <cjk>
	0xFCEF: '齩' // U+9F69 <cjk>
	0xFCF0: '𪘚' // U+2A61A <cjk>
	0xFCF1: '齭' // U+9F6D <cjk>
	0xFCF2: '齰' // U+9F70 <cjk>
	0xFCF3: '齵' // U+9F75 <cjk>
	0xFCF4: '𪚲' // U+2A6B2 <cjk>
}

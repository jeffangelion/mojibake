module mojibake

const jis_x_0213_doublebyte_0xf2 = {
	0x40: [`\u5820`].string() // U+5820 <cjk>
	0x41: [`\u5827`].string() // U+5827 <cjk>
	0x42: [`\u5832`].string() // U+5832 <cjk>
	0x43: [`\u5839`].string() // U+5839 <cjk>
	0x44: utf32_to_str(0x213C4) // U+213C4 <cjk>
	0x45: [`\u5849`].string() // U+5849 <cjk>
	0x46: [`\u584C`].string() // U+584C <cjk>
	0x47: [`\u5867`].string() // U+5867 <cjk>
	0x48: [`\u588A`].string() // U+588A <cjk>
	0x49: [`\u588B`].string() // U+588B <cjk>
	0x4A: [`\u588D`].string() // U+588D <cjk>
	0x4B: [`\u588F`].string() // U+588F <cjk>
	0x4C: [`\u5890`].string() // U+5890 <cjk>
	0x4D: [`\u5894`].string() // U+5894 <cjk>
	0x4E: [`\u589D`].string() // U+589D <cjk>
	0x4F: [`\u58AA`].string() // U+58AA <cjk>
	0x50: [`\u58B1`].string() // U+58B1 <cjk>
	0x51: utf32_to_str(0x2146D) // U+2146D <cjk>
	0x52: [`\u58C3`].string() // U+58C3 <cjk>
	0x53: [`\u58CD`].string() // U+58CD <cjk>
	0x54: [`\u58E2`].string() // U+58E2 <cjk>
	0x55: [`\u58F3`].string() // U+58F3 <cjk>
	0x56: [`\u58F4`].string() // U+58F4 <cjk>
	0x57: [`\u5905`].string() // U+5905 <cjk>
	0x58: [`\u5906`].string() // U+5906 <cjk>
	0x59: [`\u590B`].string() // U+590B <cjk>
	0x5A: [`\u590D`].string() // U+590D <cjk>
	0x5B: [`\u5914`].string() // U+5914 <cjk>
	0x5C: [`\u5924`].string() // U+5924 <cjk>
	0x5D: utf32_to_str(0x215D7) // U+215D7 <cjk>
	0x5E: [`\u3691`].string() // U+3691 <cjk>
	0x5F: [`\u593D`].string() // U+593D <cjk>
	0x60: [`\u3699`].string() // U+3699 <cjk>
	0x61: [`\u5946`].string() // U+5946 <cjk>
	0x62: [`\u3696`].string() // U+3696 <cjk>
	0x63: utf32_to_str(0x26C29) // U+26C29 <cjk>
	0x64: [`\u595B`].string() // U+595B <cjk>
	0x65: [`\u595F`].string() // U+595F <cjk>
	0x66: utf32_to_str(0x21647) // U+21647 <cjk>
	0x67: [`\u5975`].string() // U+5975 <cjk>
	0x68: [`\u5976`].string() // U+5976 <cjk>
	0x69: [`\u597C`].string() // U+597C <cjk>
	0x6A: [`\u599F`].string() // U+599F <cjk>
	0x6B: [`\u59AE`].string() // U+59AE <cjk>
	0x6C: [`\u59BC`].string() // U+59BC <cjk>
	0x6D: [`\u59C8`].string() // U+59C8 <cjk>
	0x6E: [`\u59CD`].string() // U+59CD <cjk>
	0x6F: [`\u59DE`].string() // U+59DE <cjk>
	0x70: [`\u59E3`].string() // U+59E3 <cjk>
	0x71: [`\u59E4`].string() // U+59E4 <cjk>
	0x72: [`\u59E7`].string() // U+59E7 <cjk>
	0x73: [`\u59EE`].string() // U+59EE <cjk>
	0x74: utf32_to_str(0x21706) // U+21706 <cjk>
	0x75: utf32_to_str(0x21742) // U+21742 <cjk>
	0x76: [`\u36CF`].string() // U+36CF <cjk>
	0x77: [`\u5A0C`].string() // U+5A0C <cjk>
	0x78: [`\u5A0D`].string() // U+5A0D <cjk>
	0x79: [`\u5A17`].string() // U+5A17 <cjk>
	0x7A: [`\u5A27`].string() // U+5A27 <cjk>
	0x7B: [`\u5A2D`].string() // U+5A2D <cjk>
	0x7C: [`\u5A55`].string() // U+5A55 <cjk>
	0x7D: [`\u5A65`].string() // U+5A65 <cjk>
	0x7E: [`\u5A7A`].string() // U+5A7A <cjk>
	0x80: [`\u5A8B`].string() // U+5A8B <cjk>
	0x81: [`\u5A9C`].string() // U+5A9C <cjk>
	0x82: [`\u5A9F`].string() // U+5A9F <cjk>
	0x83: [`\u5AA0`].string() // U+5AA0 <cjk>
	0x84: [`\u5AA2`].string() // U+5AA2 <cjk>
	0x85: [`\u5AB1`].string() // U+5AB1 <cjk>
	0x86: [`\u5AB3`].string() // U+5AB3 <cjk>
	0x87: [`\u5AB5`].string() // U+5AB5 <cjk>
	0x88: [`\u5ABA`].string() // U+5ABA <cjk>
	0x89: [`\u5ABF`].string() // U+5ABF <cjk>
	0x8A: [`\u5ADA`].string() // U+5ADA <cjk>
	0x8B: [`\u5ADC`].string() // U+5ADC <cjk>
	0x8C: [`\u5AE0`].string() // U+5AE0 <cjk>
	0x8D: [`\u5AE5`].string() // U+5AE5 <cjk>
	0x8E: [`\u5AF0`].string() // U+5AF0 <cjk>
	0x8F: [`\u5AEE`].string() // U+5AEE <cjk>
	0x90: [`\u5AF5`].string() // U+5AF5 <cjk>
	0x91: [`\u5B00`].string() // U+5B00 <cjk>
	0x92: [`\u5B08`].string() // U+5B08 <cjk>
	0x93: [`\u5B17`].string() // U+5B17 <cjk>
	0x94: [`\u5B34`].string() // U+5B34 <cjk>
	0x95: [`\u5B2D`].string() // U+5B2D <cjk>
	0x96: [`\u5B4C`].string() // U+5B4C <cjk>
	0x97: [`\u5B52`].string() // U+5B52 <cjk>
	0x98: [`\u5B68`].string() // U+5B68 <cjk>
	0x99: [`\u5B6F`].string() // U+5B6F <cjk>
	0x9A: [`\u5B7C`].string() // U+5B7C <cjk>
	0x9B: [`\u5B7F`].string() // U+5B7F <cjk>
	0x9C: [`\u5B81`].string() // U+5B81 <cjk>
	0x9D: [`\u5B84`].string() // U+5B84 <cjk>
	0x9E: utf32_to_str(0x219C3) // U+219C3 <cjk>
	0x9F: [`\u5E6E`].string() // U+5E6E <cjk>
	0xA0: utf32_to_str(0x2217B) // U+2217B <cjk>
	0xA1: [`\u5EA5`].string() // U+5EA5 <cjk>
	0xA2: [`\u5EAA`].string() // U+5EAA <cjk>
	0xA3: [`\u5EAC`].string() // U+5EAC <cjk>
	0xA4: [`\u5EB9`].string() // U+5EB9 <cjk>
	0xA5: [`\u5EBF`].string() // U+5EBF <cjk>
	0xA6: [`\u5EC6`].string() // U+5EC6 <cjk>
	0xA7: [`\u5ED2`].string() // U+5ED2 <cjk>
	0xA8: [`\u5ED9`].string() // U+5ED9 <cjk>
	0xA9: utf32_to_str(0x2231E) // U+2231E <cjk>
	0xAA: [`\u5EFD`].string() // U+5EFD <cjk>
	0xAB: [`\u5F08`].string() // U+5F08 <cjk>
	0xAC: [`\u5F0E`].string() // U+5F0E <cjk>
	0xAD: [`\u5F1C`].string() // U+5F1C <cjk>
	0xAE: utf32_to_str(0x223AD) // U+223AD <cjk>
	0xAF: [`\u5F1E`].string() // U+5F1E <cjk>
	0xB0: [`\u5F47`].string() // U+5F47 <cjk>
	0xB1: [`\u5F63`].string() // U+5F63 <cjk>
	0xB2: [`\u5F72`].string() // U+5F72 <cjk>
	0xB3: [`\u5F7E`].string() // U+5F7E <cjk>
	0xB4: [`\u5F8F`].string() // U+5F8F <cjk>
	0xB5: [`\u5FA2`].string() // U+5FA2 <cjk>
	0xB6: [`\u5FA4`].string() // U+5FA4 <cjk>
	0xB7: [`\u5FB8`].string() // U+5FB8 <cjk>
	0xB8: [`\u5FC4`].string() // U+5FC4 <cjk>
	0xB9: [`\u38FA`].string() // U+38FA <cjk>
	0xBA: [`\u5FC7`].string() // U+5FC7 <cjk>
	0xBB: [`\u5FCB`].string() // U+5FCB <cjk>
	0xBC: [`\u5FD2`].string() // U+5FD2 <cjk>
	0xBD: [`\u5FD3`].string() // U+5FD3 <cjk>
	0xBE: [`\u5FD4`].string() // U+5FD4 <cjk>
	0xBF: [`\u5FE2`].string() // U+5FE2 <cjk>
	0xC0: [`\u5FEE`].string() // U+5FEE <cjk>
	0xC1: [`\u5FEF`].string() // U+5FEF <cjk>
	0xC2: [`\u5FF3`].string() // U+5FF3 <cjk>
	0xC3: [`\u5FFC`].string() // U+5FFC <cjk>
	0xC4: [`\u3917`].string() // U+3917 <cjk>
	0xC5: [`\u6017`].string() // U+6017 <cjk>
	0xC6: [`\u6022`].string() // U+6022 <cjk>
	0xC7: [`\u6024`].string() // U+6024 <cjk>
	0xC8: [`\u391A`].string() // U+391A <cjk>
	0xC9: [`\u604C`].string() // U+604C <cjk>
	0xCA: [`\u607F`].string() // U+607F <cjk>
	0xCB: [`\u608A`].string() // U+608A <cjk>
	0xCC: [`\u6095`].string() // U+6095 <cjk>
	0xCD: [`\u60A8`].string() // U+60A8 <cjk>
	0xCE: utf32_to_str(0x226F3) // U+226F3 <cjk>
	0xCF: [`\u60B0`].string() // U+60B0 <cjk>
	0xD0: [`\u60B1`].string() // U+60B1 <cjk>
	0xD1: [`\u60BE`].string() // U+60BE <cjk>
	0xD2: [`\u60C8`].string() // U+60C8 <cjk>
	0xD3: [`\u60D9`].string() // U+60D9 <cjk>
	0xD4: [`\u60DB`].string() // U+60DB <cjk>
	0xD5: [`\u60EE`].string() // U+60EE <cjk>
	0xD6: [`\u60F2`].string() // U+60F2 <cjk>
	0xD7: [`\u60F5`].string() // U+60F5 <cjk>
	0xD8: [`\u6110`].string() // U+6110 <cjk>
	0xD9: [`\u6112`].string() // U+6112 <cjk>
	0xDA: [`\u6113`].string() // U+6113 <cjk>
	0xDB: [`\u6119`].string() // U+6119 <cjk>
	0xDC: [`\u611E`].string() // U+611E <cjk>
	0xDD: [`\u613A`].string() // U+613A <cjk>
	0xDE: [`\u396F`].string() // U+396F <cjk>
	0xDF: [`\u6141`].string() // U+6141 <cjk>
	0xE0: [`\u6146`].string() // U+6146 <cjk>
	0xE1: [`\u6160`].string() // U+6160 <cjk>
	0xE2: [`\u617C`].string() // U+617C <cjk>
	0xE3: utf32_to_str(0x2285B) // U+2285B <cjk>
	0xE4: [`\u6192`].string() // U+6192 <cjk>
	0xE5: [`\u6193`].string() // U+6193 <cjk>
	0xE6: [`\u6197`].string() // U+6197 <cjk>
	0xE7: [`\u6198`].string() // U+6198 <cjk>
	0xE8: [`\u61A5`].string() // U+61A5 <cjk>
	0xE9: [`\u61A8`].string() // U+61A8 <cjk>
	0xEA: [`\u61AD`].string() // U+61AD <cjk>
	0xEB: utf32_to_str(0x228AB) // U+228AB <cjk>
	0xEC: [`\u61D5`].string() // U+61D5 <cjk>
	0xED: [`\u61DD`].string() // U+61DD <cjk>
	0xEE: [`\u61DF`].string() // U+61DF <cjk>
	0xEF: [`\u61F5`].string() // U+61F5 <cjk>
	0xF0: utf32_to_str(0x2298F) // U+2298F <cjk>
	0xF1: [`\u6215`].string() // U+6215 <cjk>
	0xF2: [`\u6223`].string() // U+6223 <cjk>
	0xF3: [`\u6229`].string() // U+6229 <cjk>
	0xF4: [`\u6246`].string() // U+6246 <cjk>
	0xF5: [`\u624C`].string() // U+624C <cjk>
	0xF6: [`\u6251`].string() // U+6251 <cjk>
	0xF7: [`\u6252`].string() // U+6252 <cjk>
	0xF8: [`\u6261`].string() // U+6261 <cjk>
	0xF9: [`\u6264`].string() // U+6264 <cjk>
	0xFA: [`\u627B`].string() // U+627B <cjk>
	0xFB: [`\u626D`].string() // U+626D <cjk>
	0xFC: [`\u6273`].string() // U+6273 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x88 = {
	0x40: [`\u54A9`].string() // U+54A9 <cjk>
	0x41: [`\u54C6`].string() // U+54C6 <cjk>
	0x42: [`\u54FF`].string() // U+54FF <cjk>
	0x43: [`\u550E`].string() // U+550E <cjk>
	0x44: [`\u552B`].string() // U+552B <cjk>
	0x45: [`\u5535`].string() // U+5535 <cjk>
	0x46: [`\u5550`].string() // U+5550 <cjk>
	0x47: [`\u555E`].string() // U+555E <cjk>
	0x48: [`\u5581`].string() // U+5581 <cjk>
	0x49: [`\u5586`].string() // U+5586 <cjk>
	0x4A: [`\u558E`].string() // U+558E <cjk>
	0x4B: [`\uFA36`].string() // U+FA36 CJK COMPATIBILITY IDEOGRAPH-FA36
	0x4C: [`\u55AD`].string() // U+55AD <cjk>
	0x4D: [`\u55CE`].string() // U+55CE <cjk>
	0x4E: [`\uFA37`].string() // U+FA37 CJK COMPATIBILITY IDEOGRAPH-FA37
	0x4F: [`\u5608`].string() // U+5608 <cjk>
	0x50: [`\u560E`].string() // U+560E <cjk>
	0x51: [`\u563B`].string() // U+563B <cjk>
	0x52: [`\u5649`].string() // U+5649 <cjk>
	0x53: [`\u5676`].string() // U+5676 <cjk>
	0x54: [`\u5666`].string() // U+5666 <cjk>
	0x55: [`\uFA38`].string() // U+FA38 CJK COMPATIBILITY IDEOGRAPH-FA38
	0x56: [`\u566F`].string() // U+566F <cjk>
	0x57: [`\u5671`].string() // U+5671 <cjk>
	0x58: [`\u5672`].string() // U+5672 <cjk>
	0x59: [`\u5699`].string() // U+5699 <cjk>
	0x5A: [`\u569E`].string() // U+569E <cjk>
	0x5B: [`\u56A9`].string() // U+56A9 <cjk>
	0x5C: [`\u56AC`].string() // U+56AC <cjk>
	0x5D: [`\u56B3`].string() // U+56B3 <cjk>
	0x5E: [`\u56C9`].string() // U+56C9 <cjk>
	0x5F: [`\u56CA`].string() // U+56CA <cjk>
	0x60: [`\u570A`].string() // U+570A <cjk>
	0x61: utf32_to_str(0x2123D) // U+2123D <cjk>
	0x62: [`\u5721`].string() // U+5721 <cjk>
	0x63: [`\u572F`].string() // U+572F <cjk>
	0x64: [`\u5733`].string() // U+5733 <cjk>
	0x65: [`\u5734`].string() // U+5734 <cjk>
	0x66: [`\u5770`].string() // U+5770 <cjk>
	0x67: [`\u5777`].string() // U+5777 <cjk>
	0x68: [`\u577C`].string() // U+577C <cjk>
	0x69: [`\u579C`].string() // U+579C <cjk>
	0x6A: [`\uFA0F`].string() // U+FA0F CJK COMPATIBILITY IDEOGRAPH-FA0F
	0x6B: utf32_to_str(0x2131B) // U+2131B <cjk>
	0x6C: [`\u57B8`].string() // U+57B8 <cjk>
	0x6D: [`\u57C7`].string() // U+57C7 <cjk>
	0x6E: [`\u57C8`].string() // U+57C8 <cjk>
	0x6F: [`\u57CF`].string() // U+57CF <cjk>
	0x70: [`\u57E4`].string() // U+57E4 <cjk>
	0x71: [`\u57ED`].string() // U+57ED <cjk>
	0x72: [`\u57F5`].string() // U+57F5 <cjk>
	0x73: [`\u57F6`].string() // U+57F6 <cjk>
	0x74: [`\u57FF`].string() // U+57FF <cjk>
	0x75: [`\u5809`].string() // U+5809 <cjk>
	0x76: [`\uFA10`].string() // U+FA10 CJK COMPATIBILITY IDEOGRAPH-FA10
	0x77: [`\u5861`].string() // U+5861 <cjk>
	0x78: [`\u5864`].string() // U+5864 <cjk>
	0x79: [`\uFA39`].string() // U+FA39 CJK COMPATIBILITY IDEOGRAPH-FA39
	0x7A: [`\u587C`].string() // U+587C <cjk>
	0x7B: [`\u5889`].string() // U+5889 <cjk>
	0x7C: [`\u589E`].string() // U+589E <cjk>
	0x7D: [`\uFA3A`].string() // U+FA3A CJK COMPATIBILITY IDEOGRAPH-FA3A
	0x7E: [`\u58A9`].string() // U+58A9 <cjk>
	0x80: utf32_to_str(0x2146E) // U+2146E <cjk>
	0x81: [`\u58D2`].string() // U+58D2 <cjk>
	0x82: [`\u58CE`].string() // U+58CE <cjk>
	0x83: [`\u58D4`].string() // U+58D4 <cjk>
	0x84: [`\u58DA`].string() // U+58DA <cjk>
	0x85: [`\u58E0`].string() // U+58E0 <cjk>
	0x86: [`\u58E9`].string() // U+58E9 <cjk>
	0x87: [`\u590C`].string() // U+590C <cjk>
	0x88: [`\u8641`].string() // U+8641 <cjk>
	0x89: [`\u595D`].string() // U+595D <cjk>
	0x8A: [`\u596D`].string() // U+596D <cjk>
	0x8B: [`\u598B`].string() // U+598B <cjk>
	0x8C: [`\u5992`].string() // U+5992 <cjk>
	0x8D: [`\u59A4`].string() // U+59A4 <cjk>
	0x8E: [`\u59C3`].string() // U+59C3 <cjk>
	0x8F: [`\u59D2`].string() // U+59D2 <cjk>
	0x90: [`\u59DD`].string() // U+59DD <cjk>
	0x91: [`\u5A13`].string() // U+5A13 <cjk>
	0x92: [`\u5A23`].string() // U+5A23 <cjk>
	0x93: [`\u5A67`].string() // U+5A67 <cjk>
	0x94: [`\u5A6D`].string() // U+5A6D <cjk>
	0x95: [`\u5A77`].string() // U+5A77 <cjk>
	0x96: [`\u5A7E`].string() // U+5A7E <cjk>
	0x97: [`\u5A84`].string() // U+5A84 <cjk>
	0x98: [`\u5A9E`].string() // U+5A9E <cjk>
	0x99: [`\u5AA7`].string() // U+5AA7 <cjk>
	0x9A: [`\u5AC4`].string() // U+5AC4 <cjk>
	0x9B: utf32_to_str(0x218BD) // U+218BD <cjk>
	0x9C: [`\u5B19`].string() // U+5B19 <cjk>
	0x9D: [`\u5B25`].string() // U+5B25 <cjk>
	0x9E: [`\u525D`].string() // U+525D <cjk>
	0x9F: [`\u4E9C`].string() // U+4E9C <cjk>
	0xA0: [`\u5516`].string() // U+5516 <cjk>
	0xA1: [`\u5A03`].string() // U+5A03 <cjk>
	0xA2: [`\u963F`].string() // U+963F <cjk>
	0xA3: [`\u54C0`].string() // U+54C0 <cjk>
	0xA4: [`\u611B`].string() // U+611B <cjk>
	0xA5: [`\u6328`].string() // U+6328 <cjk>
	0xA6: [`\u59F6`].string() // U+59F6 <cjk>
	0xA7: [`\u9022`].string() // U+9022 <cjk>
	0xA8: [`\u8475`].string() // U+8475 <cjk>
	0xA9: [`\u831C`].string() // U+831C <cjk>
	0xAA: [`\u7A50`].string() // U+7A50 <cjk>
	0xAB: [`\u60AA`].string() // U+60AA <cjk>
	0xAC: [`\u63E1`].string() // U+63E1 <cjk>
	0xAD: [`\u6E25`].string() // U+6E25 <cjk>
	0xAE: [`\u65ED`].string() // U+65ED <cjk>
	0xAF: [`\u8466`].string() // U+8466 <cjk>
	0xB0: [`\u82A6`].string() // U+82A6 <cjk>
	0xB1: [`\u9BF5`].string() // U+9BF5 <cjk>
	0xB2: [`\u6893`].string() // U+6893 <cjk>
	0xB3: [`\u5727`].string() // U+5727 <cjk>
	0xB4: [`\u65A1`].string() // U+65A1 <cjk>
	0xB5: [`\u6271`].string() // U+6271 <cjk>
	0xB6: [`\u5B9B`].string() // U+5B9B <cjk>
	0xB7: [`\u59D0`].string() // U+59D0 <cjk>
	0xB8: [`\u867B`].string() // U+867B <cjk>
	0xB9: [`\u98F4`].string() // U+98F4 <cjk>
	0xBA: [`\u7D62`].string() // U+7D62 <cjk>
	0xBB: [`\u7DBE`].string() // U+7DBE <cjk>
	0xBC: [`\u9B8E`].string() // U+9B8E <cjk>
	0xBD: [`\u6216`].string() // U+6216 <cjk>
	0xBE: [`\u7C9F`].string() // U+7C9F <cjk>
	0xBF: [`\u88B7`].string() // U+88B7 <cjk>
	0xC0: [`\u5B89`].string() // U+5B89 <cjk>
	0xC1: [`\u5EB5`].string() // U+5EB5 <cjk>
	0xC2: [`\u6309`].string() // U+6309 <cjk>
	0xC3: [`\u6697`].string() // U+6697 <cjk>
	0xC4: [`\u6848`].string() // U+6848 <cjk>
	0xC5: [`\u95C7`].string() // U+95C7 <cjk>
	0xC6: [`\u978D`].string() // U+978D <cjk>
	0xC7: [`\u674F`].string() // U+674F <cjk>
	0xC8: [`\u4EE5`].string() // U+4EE5 <cjk>
	0xC9: [`\u4F0A`].string() // U+4F0A <cjk>
	0xCA: [`\u4F4D`].string() // U+4F4D <cjk>
	0xCB: [`\u4F9D`].string() // U+4F9D <cjk>
	0xCC: [`\u5049`].string() // U+5049 <cjk>
	0xCD: [`\u56F2`].string() // U+56F2 <cjk>
	0xCE: [`\u5937`].string() // U+5937 <cjk>
	0xCF: [`\u59D4`].string() // U+59D4 <cjk>
	0xD0: [`\u5A01`].string() // U+5A01 <cjk>
	0xD1: [`\u5C09`].string() // U+5C09 <cjk>
	0xD2: [`\u60DF`].string() // U+60DF <cjk>
	0xD3: [`\u610F`].string() // U+610F <cjk>
	0xD4: [`\u6170`].string() // U+6170 <cjk>
	0xD5: [`\u6613`].string() // U+6613 <cjk>
	0xD6: [`\u6905`].string() // U+6905 <cjk>
	0xD7: [`\u70BA`].string() // U+70BA <cjk>
	0xD8: [`\u754F`].string() // U+754F <cjk>
	0xD9: [`\u7570`].string() // U+7570 <cjk>
	0xDA: [`\u79FB`].string() // U+79FB <cjk>
	0xDB: [`\u7DAD`].string() // U+7DAD <cjk>
	0xDC: [`\u7DEF`].string() // U+7DEF <cjk>
	0xDD: [`\u80C3`].string() // U+80C3 <cjk>
	0xDE: [`\u840E`].string() // U+840E <cjk>
	0xDF: [`\u8863`].string() // U+8863 <cjk>
	0xE0: [`\u8B02`].string() // U+8B02 <cjk>
	0xE1: [`\u9055`].string() // U+9055 <cjk>
	0xE2: [`\u907A`].string() // U+907A <cjk>
	0xE3: [`\u533B`].string() // U+533B <cjk>
	0xE4: [`\u4E95`].string() // U+4E95 <cjk>
	0xE5: [`\u4EA5`].string() // U+4EA5 <cjk>
	0xE6: [`\u57DF`].string() // U+57DF <cjk>
	0xE7: [`\u80B2`].string() // U+80B2 <cjk>
	0xE8: [`\u90C1`].string() // U+90C1 <cjk>
	0xE9: [`\u78EF`].string() // U+78EF <cjk>
	0xEA: [`\u4E00`].string() // U+4E00 <cjk>
	0xEB: [`\u58F1`].string() // U+58F1 <cjk>
	0xEC: [`\u6EA2`].string() // U+6EA2 <cjk>
	0xED: [`\u9038`].string() // U+9038 <cjk>
	0xEE: [`\u7A32`].string() // U+7A32 <cjk>
	0xEF: [`\u8328`].string() // U+8328 <cjk>
	0xF0: [`\u828B`].string() // U+828B <cjk>
	0xF1: [`\u9C2F`].string() // U+9C2F <cjk>
	0xF2: [`\u5141`].string() // U+5141 <cjk>
	0xF3: [`\u5370`].string() // U+5370 <cjk>
	0xF4: [`\u54BD`].string() // U+54BD <cjk>
	0xF5: [`\u54E1`].string() // U+54E1 <cjk>
	0xF6: [`\u56E0`].string() // U+56E0 <cjk>
	0xF7: [`\u59FB`].string() // U+59FB <cjk>
	0xF8: [`\u5F15`].string() // U+5F15 <cjk>
	0xF9: [`\u98F2`].string() // U+98F2 <cjk>
	0xFA: [`\u6DEB`].string() // U+6DEB <cjk>
	0xFB: [`\u80E4`].string() // U+80E4 <cjk>
	0xFC: [`\u852D`].string() // U+852D <cjk>
}

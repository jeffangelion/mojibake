module mojibake

const jis_x_0213_doublebyte_0x9f = {
	0x40: [`\u6A97`].string() // U+6A97 <cjk>
	0x41: [`\u8617`].string() // U+8617 <cjk>
	0x42: [`\u6ABB`].string() // U+6ABB <cjk>
	0x43: [`\u6AC3`].string() // U+6AC3 <cjk>
	0x44: [`\u6AC2`].string() // U+6AC2 <cjk>
	0x45: [`\u6AB8`].string() // U+6AB8 <cjk>
	0x46: [`\u6AB3`].string() // U+6AB3 <cjk>
	0x47: [`\u6AAC`].string() // U+6AAC <cjk>
	0x48: [`\u6ADE`].string() // U+6ADE <cjk>
	0x49: [`\u6AD1`].string() // U+6AD1 <cjk>
	0x4A: [`\u6ADF`].string() // U+6ADF <cjk>
	0x4B: [`\u6AAA`].string() // U+6AAA <cjk>
	0x4C: [`\u6ADA`].string() // U+6ADA <cjk>
	0x4D: [`\u6AEA`].string() // U+6AEA <cjk>
	0x4E: [`\u6AFB`].string() // U+6AFB <cjk>
	0x4F: [`\u6B05`].string() // U+6B05 <cjk>
	0x50: [`\u8616`].string() // U+8616 <cjk>
	0x51: [`\u6AFA`].string() // U+6AFA <cjk>
	0x52: [`\u6B12`].string() // U+6B12 <cjk>
	0x53: [`\u6B16`].string() // U+6B16 <cjk>
	0x54: [`\u9B31`].string() // U+9B31 <cjk>
	0x55: [`\u6B1F`].string() // U+6B1F <cjk>
	0x56: [`\u6B38`].string() // U+6B38 <cjk>
	0x57: [`\u6B37`].string() // U+6B37 <cjk>
	0x58: [`\u76DC`].string() // U+76DC <cjk>
	0x59: [`\u6B39`].string() // U+6B39 <cjk>
	0x5A: [`\u98EE`].string() // U+98EE <cjk>
	0x5B: [`\u6B47`].string() // U+6B47 <cjk>
	0x5C: [`\u6B43`].string() // U+6B43 <cjk>
	0x5D: [`\u6B49`].string() // U+6B49 <cjk>
	0x5E: [`\u6B50`].string() // U+6B50 <cjk>
	0x5F: [`\u6B59`].string() // U+6B59 <cjk>
	0x60: [`\u6B54`].string() // U+6B54 <cjk>
	0x61: [`\u6B5B`].string() // U+6B5B <cjk>
	0x62: [`\u6B5F`].string() // U+6B5F <cjk>
	0x63: [`\u6B61`].string() // U+6B61 <cjk>
	0x64: [`\u6B78`].string() // U+6B78 <cjk>
	0x65: [`\u6B79`].string() // U+6B79 <cjk>
	0x66: [`\u6B7F`].string() // U+6B7F <cjk>
	0x67: [`\u6B80`].string() // U+6B80 <cjk>
	0x68: [`\u6B84`].string() // U+6B84 <cjk>
	0x69: [`\u6B83`].string() // U+6B83 <cjk>
	0x6A: [`\u6B8D`].string() // U+6B8D <cjk>
	0x6B: [`\u6B98`].string() // U+6B98 <cjk>
	0x6C: [`\u6B95`].string() // U+6B95 <cjk>
	0x6D: [`\u6B9E`].string() // U+6B9E <cjk>
	0x6E: [`\u6BA4`].string() // U+6BA4 <cjk>
	0x6F: [`\u6BAA`].string() // U+6BAA <cjk>
	0x70: [`\u6BAB`].string() // U+6BAB <cjk>
	0x71: [`\u6BAF`].string() // U+6BAF <cjk>
	0x72: [`\u6BB2`].string() // U+6BB2 <cjk>
	0x73: [`\u6BB1`].string() // U+6BB1 <cjk>
	0x74: [`\u6BB3`].string() // U+6BB3 <cjk>
	0x75: [`\u6BB7`].string() // U+6BB7 <cjk>
	0x76: [`\u6BBC`].string() // U+6BBC <cjk>
	0x77: [`\u6BC6`].string() // U+6BC6 <cjk>
	0x78: [`\u6BCB`].string() // U+6BCB <cjk>
	0x79: [`\u6BD3`].string() // U+6BD3 <cjk>
	0x7A: [`\u6BDF`].string() // U+6BDF <cjk>
	0x7B: [`\u6BEC`].string() // U+6BEC <cjk>
	0x7C: [`\u6BEB`].string() // U+6BEB <cjk>
	0x7D: [`\u6BF3`].string() // U+6BF3 <cjk>
	0x7E: [`\u6BEF`].string() // U+6BEF <cjk>
	0x80: [`\u9EBE`].string() // U+9EBE <cjk>
	0x81: [`\u6C08`].string() // U+6C08 <cjk>
	0x82: [`\u6C13`].string() // U+6C13 <cjk>
	0x83: [`\u6C14`].string() // U+6C14 <cjk>
	0x84: [`\u6C1B`].string() // U+6C1B <cjk>
	0x85: [`\u6C24`].string() // U+6C24 <cjk>
	0x86: [`\u6C23`].string() // U+6C23 <cjk>
	0x87: [`\u6C5E`].string() // U+6C5E <cjk>
	0x88: [`\u6C55`].string() // U+6C55 <cjk>
	0x89: [`\u6C62`].string() // U+6C62 <cjk>
	0x8A: [`\u6C6A`].string() // U+6C6A <cjk>
	0x8B: [`\u6C82`].string() // U+6C82 <cjk>
	0x8C: [`\u6C8D`].string() // U+6C8D <cjk>
	0x8D: [`\u6C9A`].string() // U+6C9A <cjk>
	0x8E: [`\u6C81`].string() // U+6C81 <cjk>
	0x8F: [`\u6C9B`].string() // U+6C9B <cjk>
	0x90: [`\u6C7E`].string() // U+6C7E <cjk>
	0x91: [`\u6C68`].string() // U+6C68 <cjk>
	0x92: [`\u6C73`].string() // U+6C73 <cjk>
	0x93: [`\u6C92`].string() // U+6C92 <cjk>
	0x94: [`\u6C90`].string() // U+6C90 <cjk>
	0x95: [`\u6CC4`].string() // U+6CC4 <cjk>
	0x96: [`\u6CF1`].string() // U+6CF1 <cjk>
	0x97: [`\u6CD3`].string() // U+6CD3 <cjk>
	0x98: [`\u6CBD`].string() // U+6CBD <cjk>
	0x99: [`\u6CD7`].string() // U+6CD7 <cjk>
	0x9A: [`\u6CC5`].string() // U+6CC5 <cjk>
	0x9B: [`\u6CDD`].string() // U+6CDD <cjk>
	0x9C: [`\u6CAE`].string() // U+6CAE <cjk>
	0x9D: [`\u6CB1`].string() // U+6CB1 <cjk>
	0x9E: [`\u6CBE`].string() // U+6CBE <cjk>
	0x9F: [`\u6CBA`].string() // U+6CBA <cjk>
	0xA0: [`\u6CDB`].string() // U+6CDB <cjk>
	0xA1: [`\u6CEF`].string() // U+6CEF <cjk>
	0xA2: [`\u6CD9`].string() // U+6CD9 <cjk>
	0xA3: [`\u6CEA`].string() // U+6CEA <cjk>
	0xA4: [`\u6D1F`].string() // U+6D1F <cjk>
	0xA5: [`\u884D`].string() // U+884D <cjk>
	0xA6: [`\u6D36`].string() // U+6D36 <cjk>
	0xA7: [`\u6D2B`].string() // U+6D2B <cjk>
	0xA8: [`\u6D3D`].string() // U+6D3D <cjk>
	0xA9: [`\u6D38`].string() // U+6D38 <cjk>
	0xAA: [`\u6D19`].string() // U+6D19 <cjk>
	0xAB: [`\u6D35`].string() // U+6D35 <cjk>
	0xAC: [`\u6D33`].string() // U+6D33 <cjk>
	0xAD: [`\u6D12`].string() // U+6D12 <cjk>
	0xAE: [`\u6D0C`].string() // U+6D0C <cjk>
	0xAF: [`\u6D63`].string() // U+6D63 <cjk>
	0xB0: [`\u6D93`].string() // U+6D93 <cjk>
	0xB1: [`\u6D64`].string() // U+6D64 <cjk>
	0xB2: [`\u6D5A`].string() // U+6D5A <cjk>
	0xB3: [`\u6D79`].string() // U+6D79 <cjk>
	0xB4: [`\u6D59`].string() // U+6D59 <cjk>
	0xB5: [`\u6D8E`].string() // U+6D8E <cjk>
	0xB6: [`\u6D95`].string() // U+6D95 <cjk>
	0xB7: [`\u6FE4`].string() // U+6FE4 <cjk>
	0xB8: [`\u6D85`].string() // U+6D85 <cjk>
	0xB9: [`\u6DF9`].string() // U+6DF9 <cjk>
	0xBA: [`\u6E15`].string() // U+6E15 <cjk>
	0xBB: [`\u6E0A`].string() // U+6E0A <cjk>
	0xBC: [`\u6DB5`].string() // U+6DB5 <cjk>
	0xBD: [`\u6DC7`].string() // U+6DC7 <cjk>
	0xBE: [`\u6DE6`].string() // U+6DE6 <cjk>
	0xBF: [`\u6DB8`].string() // U+6DB8 <cjk>
	0xC0: [`\u6DC6`].string() // U+6DC6 <cjk>
	0xC1: [`\u6DEC`].string() // U+6DEC <cjk>
	0xC2: [`\u6DDE`].string() // U+6DDE <cjk>
	0xC3: [`\u6DCC`].string() // U+6DCC <cjk>
	0xC4: [`\u6DE8`].string() // U+6DE8 <cjk>
	0xC5: [`\u6DD2`].string() // U+6DD2 <cjk>
	0xC6: [`\u6DC5`].string() // U+6DC5 <cjk>
	0xC7: [`\u6DFA`].string() // U+6DFA <cjk>
	0xC8: [`\u6DD9`].string() // U+6DD9 <cjk>
	0xC9: [`\u6DE4`].string() // U+6DE4 <cjk>
	0xCA: [`\u6DD5`].string() // U+6DD5 <cjk>
	0xCB: [`\u6DEA`].string() // U+6DEA <cjk>
	0xCC: [`\u6DEE`].string() // U+6DEE <cjk>
	0xCD: [`\u6E2D`].string() // U+6E2D <cjk>
	0xCE: [`\u6E6E`].string() // U+6E6E <cjk>
	0xCF: [`\u6E2E`].string() // U+6E2E <cjk>
	0xD0: [`\u6E19`].string() // U+6E19 <cjk>
	0xD1: [`\u6E72`].string() // U+6E72 <cjk>
	0xD2: [`\u6E5F`].string() // U+6E5F <cjk>
	0xD3: [`\u6E3E`].string() // U+6E3E <cjk>
	0xD4: [`\u6E23`].string() // U+6E23 <cjk>
	0xD5: [`\u6E6B`].string() // U+6E6B <cjk>
	0xD6: [`\u6E2B`].string() // U+6E2B <cjk>
	0xD7: [`\u6E76`].string() // U+6E76 <cjk>
	0xD8: [`\u6E4D`].string() // U+6E4D <cjk>
	0xD9: [`\u6E1F`].string() // U+6E1F <cjk>
	0xDA: [`\u6E43`].string() // U+6E43 <cjk>
	0xDB: [`\u6E3A`].string() // U+6E3A <cjk>
	0xDC: [`\u6E4E`].string() // U+6E4E <cjk>
	0xDD: [`\u6E24`].string() // U+6E24 <cjk>
	0xDE: [`\u6EFF`].string() // U+6EFF <cjk>
	0xDF: [`\u6E1D`].string() // U+6E1D <cjk>
	0xE0: [`\u6E38`].string() // U+6E38 <cjk>
	0xE1: [`\u6E82`].string() // U+6E82 <cjk>
	0xE2: [`\u6EAA`].string() // U+6EAA <cjk>
	0xE3: [`\u6E98`].string() // U+6E98 <cjk>
	0xE4: [`\u6EC9`].string() // U+6EC9 <cjk>
	0xE5: [`\u6EB7`].string() // U+6EB7 <cjk>
	0xE6: [`\u6ED3`].string() // U+6ED3 <cjk>
	0xE7: [`\u6EBD`].string() // U+6EBD <cjk>
	0xE8: [`\u6EAF`].string() // U+6EAF <cjk>
	0xE9: [`\u6EC4`].string() // U+6EC4 <cjk>
	0xEA: [`\u6EB2`].string() // U+6EB2 <cjk>
	0xEB: [`\u6ED4`].string() // U+6ED4 <cjk>
	0xEC: [`\u6ED5`].string() // U+6ED5 <cjk>
	0xED: [`\u6E8F`].string() // U+6E8F <cjk>
	0xEE: [`\u6EA5`].string() // U+6EA5 <cjk>
	0xEF: [`\u6EC2`].string() // U+6EC2 <cjk>
	0xF0: [`\u6E9F`].string() // U+6E9F <cjk>
	0xF1: [`\u6F41`].string() // U+6F41 <cjk>
	0xF2: [`\u6F11`].string() // U+6F11 <cjk>
	0xF3: [`\u704C`].string() // U+704C <cjk>
	0xF4: [`\u6EEC`].string() // U+6EEC <cjk>
	0xF5: [`\u6EF8`].string() // U+6EF8 <cjk>
	0xF6: [`\u6EFE`].string() // U+6EFE <cjk>
	0xF7: [`\u6F3F`].string() // U+6F3F <cjk>
	0xF8: [`\u6EF2`].string() // U+6EF2 <cjk>
	0xF9: [`\u6F31`].string() // U+6F31 <cjk>
	0xFA: [`\u6EEF`].string() // U+6EEF <cjk>
	0xFB: [`\u6F32`].string() // U+6F32 <cjk>
	0xFC: [`\u6ECC`].string() // U+6ECC <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xe3 = {
	0x40: [`\u7D02`].string() // U+7D02 <cjk>
	0x41: [`\u7D1C`].string() // U+7D1C <cjk>
	0x42: [`\u7D15`].string() // U+7D15 <cjk>
	0x43: [`\u7D0A`].string() // U+7D0A <cjk>
	0x44: [`\u7D45`].string() // U+7D45 <cjk>
	0x45: [`\u7D4B`].string() // U+7D4B <cjk>
	0x46: [`\u7D2E`].string() // U+7D2E <cjk>
	0x47: [`\u7D32`].string() // U+7D32 <cjk>
	0x48: [`\u7D3F`].string() // U+7D3F <cjk>
	0x49: [`\u7D35`].string() // U+7D35 <cjk>
	0x4A: [`\u7D46`].string() // U+7D46 <cjk>
	0x4B: [`\u7D73`].string() // U+7D73 <cjk>
	0x4C: [`\u7D56`].string() // U+7D56 <cjk>
	0x4D: [`\u7D4E`].string() // U+7D4E <cjk>
	0x4E: [`\u7D72`].string() // U+7D72 <cjk>
	0x4F: [`\u7D68`].string() // U+7D68 <cjk>
	0x50: [`\u7D6E`].string() // U+7D6E <cjk>
	0x51: [`\u7D4F`].string() // U+7D4F <cjk>
	0x52: [`\u7D63`].string() // U+7D63 <cjk>
	0x53: [`\u7D93`].string() // U+7D93 <cjk>
	0x54: [`\u7D89`].string() // U+7D89 <cjk>
	0x55: [`\u7D5B`].string() // U+7D5B <cjk>
	0x56: [`\u7D8F`].string() // U+7D8F <cjk>
	0x57: [`\u7D7D`].string() // U+7D7D <cjk>
	0x58: [`\u7D9B`].string() // U+7D9B <cjk>
	0x59: [`\u7DBA`].string() // U+7DBA <cjk>
	0x5A: [`\u7DAE`].string() // U+7DAE <cjk>
	0x5B: [`\u7DA3`].string() // U+7DA3 <cjk>
	0x5C: [`\u7DB5`].string() // U+7DB5 <cjk>
	0x5D: [`\u7DC7`].string() // U+7DC7 <cjk>
	0x5E: [`\u7DBD`].string() // U+7DBD <cjk>
	0x5F: [`\u7DAB`].string() // U+7DAB <cjk>
	0x60: [`\u7E3D`].string() // U+7E3D <cjk>
	0x61: [`\u7DA2`].string() // U+7DA2 <cjk>
	0x62: [`\u7DAF`].string() // U+7DAF <cjk>
	0x63: [`\u7DDC`].string() // U+7DDC <cjk>
	0x64: [`\u7DB8`].string() // U+7DB8 <cjk>
	0x65: [`\u7D9F`].string() // U+7D9F <cjk>
	0x66: [`\u7DB0`].string() // U+7DB0 <cjk>
	0x67: [`\u7DD8`].string() // U+7DD8 <cjk>
	0x68: [`\u7DDD`].string() // U+7DDD <cjk>
	0x69: [`\u7DE4`].string() // U+7DE4 <cjk>
	0x6A: [`\u7DDE`].string() // U+7DDE <cjk>
	0x6B: [`\u7DFB`].string() // U+7DFB <cjk>
	0x6C: [`\u7DF2`].string() // U+7DF2 <cjk>
	0x6D: [`\u7DE1`].string() // U+7DE1 <cjk>
	0x6E: [`\u7E05`].string() // U+7E05 <cjk>
	0x6F: [`\u7E0A`].string() // U+7E0A <cjk>
	0x70: [`\u7E23`].string() // U+7E23 <cjk>
	0x71: [`\u7E21`].string() // U+7E21 <cjk>
	0x72: [`\u7E12`].string() // U+7E12 <cjk>
	0x73: [`\u7E31`].string() // U+7E31 <cjk>
	0x74: [`\u7E1F`].string() // U+7E1F <cjk>
	0x75: [`\u7E09`].string() // U+7E09 <cjk>
	0x76: [`\u7E0B`].string() // U+7E0B <cjk>
	0x77: [`\u7E22`].string() // U+7E22 <cjk>
	0x78: [`\u7E46`].string() // U+7E46 <cjk>
	0x79: [`\u7E66`].string() // U+7E66 <cjk>
	0x7A: [`\u7E3B`].string() // U+7E3B <cjk>
	0x7B: [`\u7E35`].string() // U+7E35 <cjk>
	0x7C: [`\u7E39`].string() // U+7E39 <cjk>
	0x7D: [`\u7E43`].string() // U+7E43 <cjk>
	0x7E: [`\u7E37`].string() // U+7E37 <cjk>
	0x80: [`\u7E32`].string() // U+7E32 <cjk>
	0x81: [`\u7E3A`].string() // U+7E3A <cjk>
	0x82: [`\u7E67`].string() // U+7E67 <cjk>
	0x83: [`\u7E5D`].string() // U+7E5D <cjk>
	0x84: [`\u7E56`].string() // U+7E56 <cjk>
	0x85: [`\u7E5E`].string() // U+7E5E <cjk>
	0x86: [`\u7E59`].string() // U+7E59 <cjk>
	0x87: [`\u7E5A`].string() // U+7E5A <cjk>
	0x88: [`\u7E79`].string() // U+7E79 <cjk>
	0x89: [`\u7E6A`].string() // U+7E6A <cjk>
	0x8A: [`\u7E69`].string() // U+7E69 <cjk>
	0x8B: [`\u7E7C`].string() // U+7E7C <cjk>
	0x8C: [`\u7E7B`].string() // U+7E7B <cjk>
	0x8D: [`\u7E83`].string() // U+7E83 <cjk>
	0x8E: [`\u7DD5`].string() // U+7DD5 <cjk>
	0x8F: [`\u7E7D`].string() // U+7E7D <cjk>
	0x90: [`\u8FAE`].string() // U+8FAE <cjk>
	0x91: [`\u7E7F`].string() // U+7E7F <cjk>
	0x92: [`\u7E88`].string() // U+7E88 <cjk>
	0x93: [`\u7E89`].string() // U+7E89 <cjk>
	0x94: [`\u7E8C`].string() // U+7E8C <cjk>
	0x95: [`\u7E92`].string() // U+7E92 <cjk>
	0x96: [`\u7E90`].string() // U+7E90 <cjk>
	0x97: [`\u7E93`].string() // U+7E93 <cjk>
	0x98: [`\u7E94`].string() // U+7E94 <cjk>
	0x99: [`\u7E96`].string() // U+7E96 <cjk>
	0x9A: [`\u7E8E`].string() // U+7E8E <cjk>
	0x9B: [`\u7E9B`].string() // U+7E9B <cjk>
	0x9C: [`\u7E9C`].string() // U+7E9C <cjk>
	0x9D: [`\u7F38`].string() // U+7F38 <cjk>
	0x9E: [`\u7F3A`].string() // U+7F3A <cjk>
	0x9F: [`\u7F45`].string() // U+7F45 <cjk>
	0xA0: [`\u7F4C`].string() // U+7F4C <cjk>
	0xA1: [`\u7F4D`].string() // U+7F4D <cjk>
	0xA2: [`\u7F4E`].string() // U+7F4E <cjk>
	0xA3: [`\u7F50`].string() // U+7F50 <cjk>
	0xA4: [`\u7F51`].string() // U+7F51 <cjk>
	0xA5: [`\u7F55`].string() // U+7F55 <cjk>
	0xA6: [`\u7F54`].string() // U+7F54 <cjk>
	0xA7: [`\u7F58`].string() // U+7F58 <cjk>
	0xA8: [`\u7F5F`].string() // U+7F5F <cjk>
	0xA9: [`\u7F60`].string() // U+7F60 <cjk>
	0xAA: [`\u7F68`].string() // U+7F68 <cjk>
	0xAB: [`\u7F69`].string() // U+7F69 <cjk>
	0xAC: [`\u7F67`].string() // U+7F67 <cjk>
	0xAD: [`\u7F78`].string() // U+7F78 <cjk>
	0xAE: [`\u7F82`].string() // U+7F82 <cjk>
	0xAF: [`\u7F86`].string() // U+7F86 <cjk>
	0xB0: [`\u7F83`].string() // U+7F83 <cjk>
	0xB1: [`\u7F88`].string() // U+7F88 <cjk>
	0xB2: [`\u7F87`].string() // U+7F87 <cjk>
	0xB3: [`\u7F8C`].string() // U+7F8C <cjk>
	0xB4: [`\u7F94`].string() // U+7F94 <cjk>
	0xB5: [`\u7F9E`].string() // U+7F9E <cjk>
	0xB6: [`\u7F9D`].string() // U+7F9D <cjk>
	0xB7: [`\u7F9A`].string() // U+7F9A <cjk>
	0xB8: [`\u7FA3`].string() // U+7FA3 <cjk>
	0xB9: [`\u7FAF`].string() // U+7FAF <cjk>
	0xBA: [`\u7FB2`].string() // U+7FB2 <cjk>
	0xBB: [`\u7FB9`].string() // U+7FB9 <cjk>
	0xBC: [`\u7FAE`].string() // U+7FAE <cjk>
	0xBD: [`\u7FB6`].string() // U+7FB6 <cjk>
	0xBE: [`\u7FB8`].string() // U+7FB8 <cjk>
	0xBF: [`\u8B71`].string() // U+8B71 <cjk>
	0xC0: [`\u7FC5`].string() // U+7FC5 <cjk>
	0xC1: [`\u7FC6`].string() // U+7FC6 <cjk>
	0xC2: [`\u7FCA`].string() // U+7FCA <cjk>
	0xC3: [`\u7FD5`].string() // U+7FD5 <cjk>
	0xC4: [`\u7FD4`].string() // U+7FD4 <cjk>
	0xC5: [`\u7FE1`].string() // U+7FE1 <cjk>
	0xC6: [`\u7FE6`].string() // U+7FE6 <cjk>
	0xC7: [`\u7FE9`].string() // U+7FE9 <cjk>
	0xC8: [`\u7FF3`].string() // U+7FF3 <cjk>
	0xC9: [`\u7FF9`].string() // U+7FF9 <cjk>
	0xCA: [`\u98DC`].string() // U+98DC <cjk>
	0xCB: [`\u8006`].string() // U+8006 <cjk>
	0xCC: [`\u8004`].string() // U+8004 <cjk>
	0xCD: [`\u800B`].string() // U+800B <cjk>
	0xCE: [`\u8012`].string() // U+8012 <cjk>
	0xCF: [`\u8018`].string() // U+8018 <cjk>
	0xD0: [`\u8019`].string() // U+8019 <cjk>
	0xD1: [`\u801C`].string() // U+801C <cjk>
	0xD2: [`\u8021`].string() // U+8021 <cjk>
	0xD3: [`\u8028`].string() // U+8028 <cjk>
	0xD4: [`\u803F`].string() // U+803F <cjk>
	0xD5: [`\u803B`].string() // U+803B <cjk>
	0xD6: [`\u804A`].string() // U+804A <cjk>
	0xD7: [`\u8046`].string() // U+8046 <cjk>
	0xD8: [`\u8052`].string() // U+8052 <cjk>
	0xD9: [`\u8058`].string() // U+8058 <cjk>
	0xDA: [`\u805A`].string() // U+805A <cjk>
	0xDB: [`\u805F`].string() // U+805F <cjk>
	0xDC: [`\u8062`].string() // U+8062 <cjk>
	0xDD: [`\u8068`].string() // U+8068 <cjk>
	0xDE: [`\u8073`].string() // U+8073 <cjk>
	0xDF: [`\u8072`].string() // U+8072 <cjk>
	0xE0: [`\u8070`].string() // U+8070 <cjk>
	0xE1: [`\u8076`].string() // U+8076 <cjk>
	0xE2: [`\u8079`].string() // U+8079 <cjk>
	0xE3: [`\u807D`].string() // U+807D <cjk>
	0xE4: [`\u807F`].string() // U+807F <cjk>
	0xE5: [`\u8084`].string() // U+8084 <cjk>
	0xE6: [`\u8086`].string() // U+8086 <cjk>
	0xE7: [`\u8085`].string() // U+8085 <cjk>
	0xE8: [`\u809B`].string() // U+809B <cjk>
	0xE9: [`\u8093`].string() // U+8093 <cjk>
	0xEA: [`\u809A`].string() // U+809A <cjk>
	0xEB: [`\u80AD`].string() // U+80AD <cjk>
	0xEC: [`\u5190`].string() // U+5190 <cjk>
	0xED: [`\u80AC`].string() // U+80AC <cjk>
	0xEE: [`\u80DB`].string() // U+80DB <cjk>
	0xEF: [`\u80E5`].string() // U+80E5 <cjk>
	0xF0: [`\u80D9`].string() // U+80D9 <cjk>
	0xF1: [`\u80DD`].string() // U+80DD <cjk>
	0xF2: [`\u80C4`].string() // U+80C4 <cjk>
	0xF3: [`\u80DA`].string() // U+80DA <cjk>
	0xF4: [`\u80D6`].string() // U+80D6 <cjk>
	0xF5: [`\u8109`].string() // U+8109 <cjk>
	0xF6: [`\u80EF`].string() // U+80EF <cjk>
	0xF7: [`\u80F1`].string() // U+80F1 <cjk>
	0xF8: [`\u811B`].string() // U+811B <cjk>
	0xF9: [`\u8129`].string() // U+8129 <cjk>
	0xFA: [`\u8123`].string() // U+8123 <cjk>
	0xFB: [`\u812F`].string() // U+812F <cjk>
	0xFC: [`\u814B`].string() // U+814B <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x84 = {
	0x40: [`\u0410`].string() // U+0410 CYRILLIC CAPITAL LETTER A
	0x41: [`\u0411`].string() // U+0411 CYRILLIC CAPITAL LETTER BE
	0x42: [`\u0412`].string() // U+0412 CYRILLIC CAPITAL LETTER VE
	0x43: [`\u0413`].string() // U+0413 CYRILLIC CAPITAL LETTER GHE
	0x44: [`\u0414`].string() // U+0414 CYRILLIC CAPITAL LETTER DE
	0x45: [`\u0415`].string() // U+0415 CYRILLIC CAPITAL LETTER IE
	0x46: [`\u0401`].string() // U+0401 CYRILLIC CAPITAL LETTER IO
	0x47: [`\u0416`].string() // U+0416 CYRILLIC CAPITAL LETTER ZHE
	0x48: [`\u0417`].string() // U+0417 CYRILLIC CAPITAL LETTER ZE
	0x49: [`\u0418`].string() // U+0418 CYRILLIC CAPITAL LETTER I
	0x4A: [`\u0419`].string() // U+0419 CYRILLIC CAPITAL LETTER SHORT I
	0x4B: [`\u041A`].string() // U+041A CYRILLIC CAPITAL LETTER KA
	0x4C: [`\u041B`].string() // U+041B CYRILLIC CAPITAL LETTER EL
	0x4D: [`\u041C`].string() // U+041C CYRILLIC CAPITAL LETTER EM
	0x4E: [`\u041D`].string() // U+041D CYRILLIC CAPITAL LETTER EN
	0x4F: [`\u041E`].string() // U+041E CYRILLIC CAPITAL LETTER O
	0x50: [`\u041F`].string() // U+041F CYRILLIC CAPITAL LETTER PE
	0x51: [`\u0420`].string() // U+0420 CYRILLIC CAPITAL LETTER ER
	0x52: [`\u0421`].string() // U+0421 CYRILLIC CAPITAL LETTER ES
	0x53: [`\u0422`].string() // U+0422 CYRILLIC CAPITAL LETTER TE
	0x54: [`\u0423`].string() // U+0423 CYRILLIC CAPITAL LETTER U
	0x55: [`\u0424`].string() // U+0424 CYRILLIC CAPITAL LETTER EF
	0x56: [`\u0425`].string() // U+0425 CYRILLIC CAPITAL LETTER HA
	0x57: [`\u0426`].string() // U+0426 CYRILLIC CAPITAL LETTER TSE
	0x58: [`\u0427`].string() // U+0427 CYRILLIC CAPITAL LETTER CHE
	0x59: [`\u0428`].string() // U+0428 CYRILLIC CAPITAL LETTER SHA
	0x5A: [`\u0429`].string() // U+0429 CYRILLIC CAPITAL LETTER SHCHA
	0x5B: [`\u042A`].string() // U+042A CYRILLIC CAPITAL LETTER HARD SIGN
	0x5C: [`\u042B`].string() // U+042B CYRILLIC CAPITAL LETTER YERU
	0x5D: [`\u042C`].string() // U+042C CYRILLIC CAPITAL LETTER SOFT SIGN
	0x5E: [`\u042D`].string() // U+042D CYRILLIC CAPITAL LETTER E
	0x5F: [`\u042E`].string() // U+042E CYRILLIC CAPITAL LETTER YU
	0x60: [`\u042F`].string() // U+042F CYRILLIC CAPITAL LETTER YA
	0x61: [`\u23BE`].string() // U+23BE DENTISTRY SYMBOL LIGHT VERTICAL AND TOP RIGHT
	0x62: [`\u23BF`].string() // U+23BF DENTISTRY SYMBOL LIGHT VERTICAL AND BOTTOM RIGHT
	0x63: [`\u23C0`].string() // U+23C0 DENTISTRY SYMBOL LIGHT VERTICAL WITH CIRCLE
	0x64: [`\u23C1`].string() // U+23C1 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL WITH CIRCLE
	0x65: [`\u23C2`].string() // U+23C2 DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL WITH CIRCLE
	0x66: [`\u23C3`].string() // U+23C3 DENTISTRY SYMBOL LIGHT VERTICAL WITH TRIANGLE
	0x67: [`\u23C4`].string() // U+23C4 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL WITH TRIANGLE
	0x68: [`\u23C5`].string() // U+23C5 DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL WITH TRIANGLE
	0x69: [`\u23C6`].string() // U+23C6 DENTISTRY SYMBOL LIGHT VERTICAL AND WAVE
	0x6A: [`\u23C7`].string() // U+23C7 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL WITH WAVE
	0x6B: [`\u23C8`].string() // U+23C8 DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL WITH WAVE
	0x6C: [`\u23C9`].string() // U+23C9 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL
	0x6D: [`\u23CA`].string() // U+23CA DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL
	0x6E: [`\u23CB`].string() // U+23CB DENTISTRY SYMBOL LIGHT VERTICAL AND TOP LEFT
	0x6F: [`\u23CC`].string() // U+23CC DENTISTRY SYMBOL LIGHT VERTICAL AND BOTTOM LEFT
	0x70: [`\u0430`].string() // U+0430 CYRILLIC SMALL LETTER A
	0x71: [`\u0431`].string() // U+0431 CYRILLIC SMALL LETTER BE
	0x72: [`\u0432`].string() // U+0432 CYRILLIC SMALL LETTER VE
	0x73: [`\u0433`].string() // U+0433 CYRILLIC SMALL LETTER GHE
	0x74: [`\u0434`].string() // U+0434 CYRILLIC SMALL LETTER DE
	0x75: [`\u0435`].string() // U+0435 CYRILLIC SMALL LETTER IE
	0x76: [`\u0451`].string() // U+0451 CYRILLIC SMALL LETTER IO
	0x77: [`\u0436`].string() // U+0436 CYRILLIC SMALL LETTER ZHE
	0x78: [`\u0437`].string() // U+0437 CYRILLIC SMALL LETTER ZE
	0x79: [`\u0438`].string() // U+0438 CYRILLIC SMALL LETTER I
	0x7A: [`\u0439`].string() // U+0439 CYRILLIC SMALL LETTER SHORT I
	0x7B: [`\u043A`].string() // U+043A CYRILLIC SMALL LETTER KA
	0x7C: [`\u043B`].string() // U+043B CYRILLIC SMALL LETTER EL
	0x7D: [`\u043C`].string() // U+043C CYRILLIC SMALL LETTER EM
	0x7E: [`\u043D`].string() // U+043D CYRILLIC SMALL LETTER EN
	0x80: [`\u043E`].string() // U+043E CYRILLIC SMALL LETTER O
	0x81: [`\u043F`].string() // U+043F CYRILLIC SMALL LETTER PE
	0x82: [`\u0440`].string() // U+0440 CYRILLIC SMALL LETTER ER
	0x83: [`\u0441`].string() // U+0441 CYRILLIC SMALL LETTER ES
	0x84: [`\u0442`].string() // U+0442 CYRILLIC SMALL LETTER TE
	0x85: [`\u0443`].string() // U+0443 CYRILLIC SMALL LETTER U
	0x86: [`\u0444`].string() // U+0444 CYRILLIC SMALL LETTER EF
	0x87: [`\u0445`].string() // U+0445 CYRILLIC SMALL LETTER HA
	0x88: [`\u0446`].string() // U+0446 CYRILLIC SMALL LETTER TSE
	0x89: [`\u0447`].string() // U+0447 CYRILLIC SMALL LETTER CHE
	0x8A: [`\u0448`].string() // U+0448 CYRILLIC SMALL LETTER SHA
	0x8B: [`\u0449`].string() // U+0449 CYRILLIC SMALL LETTER SHCHA
	0x8C: [`\u044A`].string() // U+044A CYRILLIC SMALL LETTER HARD SIGN
	0x8D: [`\u044B`].string() // U+044B CYRILLIC SMALL LETTER YERU
	0x8E: [`\u044C`].string() // U+044C CYRILLIC SMALL LETTER SOFT SIGN
	0x8F: [`\u044D`].string() // U+044D CYRILLIC SMALL LETTER E
	0x90: [`\u044E`].string() // U+044E CYRILLIC SMALL LETTER YU
	0x91: [`\u044F`].string() // U+044F CYRILLIC SMALL LETTER YA
	0x92: [`\u30F7`].string() // U+30F7 KATAKANA LETTER VA
	0x93: [`\u30F8`].string() // U+30F8 KATAKANA LETTER VI
	0x94: [`\u30F9`].string() // U+30F9 KATAKANA LETTER VE
	0x95: [`\u30FA`].string() // U+30FA KATAKANA LETTER VO
	0x96: [`\u22DA`].string() // U+22DA LESS-THAN EQUAL TO OR GREATER-THAN
	0x97: [`\u22DB`].string() // U+22DB GREATER-THAN EQUAL TO OR LESS-THAN
	0x98: [`\u2153`].string() // U+2153 VULGAR FRACTION ONE THIRD
	0x99: [`\u2154`].string() // U+2154 VULGAR FRACTION TWO THIRDS
	0x9A: [`\u2155`].string() // U+2155 VULGAR FRACTION ONE FIFTH
	0x9B: [`\u2713`].string() // U+2713 CHECK MARK
	0x9C: [`\u2318`].string() // U+2318 PLACE OF INTEREST SIGN
	0x9D: [`\u2423`].string() // U+2423 OPEN BOX
	0x9E: [`\u23CE`].string() // U+23CE RETURN SYMBOL
	0x9F: [`\u2500`].string() // U+2500 BOX DRAWINGS LIGHT HORIZONTAL
	0xA0: [`\u2502`].string() // U+2502 BOX DRAWINGS LIGHT VERTICAL
	0xA1: [`\u250C`].string() // U+250C BOX DRAWINGS LIGHT DOWN AND RIGHT
	0xA2: [`\u2510`].string() // U+2510 BOX DRAWINGS LIGHT DOWN AND LEFT
	0xA3: [`\u2518`].string() // U+2518 BOX DRAWINGS LIGHT UP AND LEFT
	0xA4: [`\u2514`].string() // U+2514 BOX DRAWINGS LIGHT UP AND RIGHT
	0xA5: [`\u251C`].string() // U+251C BOX DRAWINGS LIGHT VERTICAL AND RIGHT
	0xA6: [`\u252C`].string() // U+252C BOX DRAWINGS LIGHT DOWN AND HORIZONTAL
	0xA7: [`\u2524`].string() // U+2524 BOX DRAWINGS LIGHT VERTICAL AND LEFT
	0xA8: [`\u2534`].string() // U+2534 BOX DRAWINGS LIGHT UP AND HORIZONTAL
	0xA9: [`\u253C`].string() // U+253C BOX DRAWINGS LIGHT VERTICAL AND HORIZONTAL
	0xAA: [`\u2501`].string() // U+2501 BOX DRAWINGS HEAVY HORIZONTAL
	0xAB: [`\u2503`].string() // U+2503 BOX DRAWINGS HEAVY VERTICAL
	0xAC: [`\u250F`].string() // U+250F BOX DRAWINGS HEAVY DOWN AND RIGHT
	0xAD: [`\u2513`].string() // U+2513 BOX DRAWINGS HEAVY DOWN AND LEFT
	0xAE: [`\u251B`].string() // U+251B BOX DRAWINGS HEAVY UP AND LEFT
	0xAF: [`\u2517`].string() // U+2517 BOX DRAWINGS HEAVY UP AND RIGHT
	0xB0: [`\u2523`].string() // U+2523 BOX DRAWINGS HEAVY VERTICAL AND RIGHT
	0xB1: [`\u2533`].string() // U+2533 BOX DRAWINGS HEAVY DOWN AND HORIZONTAL
	0xB2: [`\u252B`].string() // U+252B BOX DRAWINGS HEAVY VERTICAL AND LEFT
	0xB3: [`\u253B`].string() // U+253B BOX DRAWINGS HEAVY UP AND HORIZONTAL
	0xB4: [`\u254B`].string() // U+254B BOX DRAWINGS HEAVY VERTICAL AND HORIZONTAL
	0xB5: [`\u2520`].string() // U+2520 BOX DRAWINGS VERTICAL HEAVY AND RIGHT LIGHT
	0xB6: [`\u252F`].string() // U+252F BOX DRAWINGS DOWN LIGHT AND HORIZONTAL HEAVY
	0xB7: [`\u2528`].string() // U+2528 BOX DRAWINGS VERTICAL HEAVY AND LEFT LIGHT
	0xB8: [`\u2537`].string() // U+2537 BOX DRAWINGS UP LIGHT AND HORIZONTAL HEAVY
	0xB9: [`\u253F`].string() // U+253F BOX DRAWINGS VERTICAL LIGHT AND HORIZONTAL HEAVY
	0xBA: [`\u251D`].string() // U+251D BOX DRAWINGS VERTICAL LIGHT AND RIGHT HEAVY
	0xBB: [`\u2530`].string() // U+2530 BOX DRAWINGS DOWN HEAVY AND HORIZONTAL LIGHT
	0xBC: [`\u2525`].string() // U+2525 BOX DRAWINGS VERTICAL LIGHT AND LEFT HEAVY
	0xBD: [`\u2538`].string() // U+2538 BOX DRAWINGS UP HEAVY AND HORIZONTAL LIGHT
	0xBE: [`\u2542`].string() // U+2542 BOX DRAWINGS VERTICAL HEAVY AND HORIZONTAL LIGHT
	0xBF: [`\u3251`].string() // U+3251 CIRCLED NUMBER TWENTY ONE
	0xC0: [`\u3252`].string() // U+3252 CIRCLED NUMBER TWENTY TWO
	0xC1: [`\u3253`].string() // U+3253 CIRCLED NUMBER TWENTY THREE
	0xC2: [`\u3254`].string() // U+3254 CIRCLED NUMBER TWENTY FOUR
	0xC3: [`\u3255`].string() // U+3255 CIRCLED NUMBER TWENTY FIVE
	0xC4: [`\u3256`].string() // U+3256 CIRCLED NUMBER TWENTY SIX
	0xC5: [`\u3257`].string() // U+3257 CIRCLED NUMBER TWENTY SEVEN
	0xC6: [`\u3258`].string() // U+3258 CIRCLED NUMBER TWENTY EIGHT
	0xC7: [`\u3259`].string() // U+3259 CIRCLED NUMBER TWENTY NINE
	0xC8: [`\u325A`].string() // U+325A CIRCLED NUMBER THIRTY
	0xC9: [`\u325B`].string() // U+325B CIRCLED NUMBER THIRTY ONE
	0xCA: [`\u325C`].string() // U+325C CIRCLED NUMBER THIRTY TWO
	0xCB: [`\u325D`].string() // U+325D CIRCLED NUMBER THIRTY THREE
	0xCC: [`\u325E`].string() // U+325E CIRCLED NUMBER THIRTY FOUR
	0xCD: [`\u325F`].string() // U+325F CIRCLED NUMBER THIRTY FIVE
	0xCE: [`\u32B1`].string() // U+32B1 CIRCLED NUMBER THIRTY SIX
	0xCF: [`\u32B2`].string() // U+32B2 CIRCLED NUMBER THIRTY SEVEN
	0xD0: [`\u32B3`].string() // U+32B3 CIRCLED NUMBER THIRTY EIGHT
	0xD1: [`\u32B4`].string() // U+32B4 CIRCLED NUMBER THIRTY NINE
	0xD2: [`\u32B5`].string() // U+32B5 CIRCLED NUMBER FORTY
	0xD3: [`\u32B6`].string() // U+32B6 CIRCLED NUMBER FORTY ONE
	0xD4: [`\u32B7`].string() // U+32B7 CIRCLED NUMBER FORTY TWO
	0xD5: [`\u32B8`].string() // U+32B8 CIRCLED NUMBER FORTY THREE
	0xD6: [`\u32B9`].string() // U+32B9 CIRCLED NUMBER FORTY FOUR
	0xD7: [`\u32BA`].string() // U+32BA CIRCLED NUMBER FORTY FIVE
	0xD8: [`\u32BB`].string() // U+32BB CIRCLED NUMBER FORTY SIX
	0xD9: [`\u32BC`].string() // U+32BC CIRCLED NUMBER FORTY SEVEN
	0xDA: [`\u32BD`].string() // U+32BD CIRCLED NUMBER FORTY EIGHT
	0xDB: [`\u32BE`].string() // U+32BE CIRCLED NUMBER FORTY NINE
	0xDC: [`\u32BF`].string() // U+32BF CIRCLED NUMBER FIFTY
	0xE5: [`\u25D0`].string() // U+25D0 CIRCLE WITH LEFT HALF BLACK
	0xE6: [`\u25D1`].string() // U+25D1 CIRCLE WITH RIGHT HALF BLACK
	0xE7: [`\u25D2`].string() // U+25D2 CIRCLE WITH LOWER HALF BLACK
	0xE8: [`\u25D3`].string() // U+25D3 CIRCLE WITH UPPER HALF BLACK
	0xE9: [`\u203C`].string() // U+203C DOUBLE EXCLAMATION MARK
	0xEA: [`\u2047`].string() // U+2047 DOUBLE QUESTION MARK
	0xEB: [`\u2048`].string() // U+2048 QUESTION EXCLAMATION MARK
	0xEC: [`\u2049`].string() // U+2049 EXCLAMATION QUESTION MARK
	0xED: [`\u01CD`].string() // U+01CD LATIN CAPITAL LETTER A WITH CARON
	0xEE: [`\u01CE`].string() // U+01CE LATIN SMALL LETTER A WITH CARON
	0xEF: [`\u01D0`].string() // U+01D0 LATIN SMALL LETTER I WITH CARON
	0xF0: [`\u1E3E`].string() // U+1E3E LATIN CAPITAL LETTER M WITH ACUTE
	0xF1: [`\u1E3F`].string() // U+1E3F LATIN SMALL LETTER M WITH ACUTE
	0xF2: [`\u01F8`].string() // U+01F8 LATIN CAPITAL LETTER N WITH GRAVE
	0xF3: [`\u01F9`].string() // U+01F9 LATIN SMALL LETTER N WITH GRAVE
	0xF4: [`\u01D1`].string() // U+01D1 LATIN CAPITAL LETTER O WITH CARON
	0xF5: [`\u01D2`].string() // U+01D2 LATIN SMALL LETTER O WITH CARON
	0xF6: [`\u01D4`].string() // U+01D4 LATIN SMALL LETTER U WITH CARON
	0xF7: [`\u01D6`].string() // U+01D6 LATIN SMALL LETTER U WITH DIAERESIS AND MACRON
	0xF8: [`\u01D8`].string() // U+01D8 LATIN SMALL LETTER U WITH DIAERESIS AND ACUTE
	0xF9: [`\u01DA`].string() // U+01DA LATIN SMALL LETTER U WITH DIAERESIS AND CARON
	0xFA: [`\u01DC`].string() // U+01DC LATIN SMALL LETTER U WITH DIAERESIS AND GRAVE
}

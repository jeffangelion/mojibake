module mojibake

const jis_x_0213_doublebyte_0x90 = {
	0x40: [`\u62ED`].string() // U+62ED <cjk>
	0x41: [`\u690D`].string() // U+690D <cjk>
	0x42: [`\u6B96`].string() // U+6B96 <cjk>
	0x43: [`\u71ED`].string() // U+71ED <cjk>
	0x44: [`\u7E54`].string() // U+7E54 <cjk>
	0x45: [`\u8077`].string() // U+8077 <cjk>
	0x46: [`\u8272`].string() // U+8272 <cjk>
	0x47: [`\u89E6`].string() // U+89E6 <cjk>
	0x48: [`\u98DF`].string() // U+98DF <cjk>
	0x49: [`\u8755`].string() // U+8755 <cjk>
	0x4A: [`\u8FB1`].string() // U+8FB1 <cjk>
	0x4B: [`\u5C3B`].string() // U+5C3B <cjk>
	0x4C: [`\u4F38`].string() // U+4F38 <cjk>
	0x4D: [`\u4FE1`].string() // U+4FE1 <cjk>
	0x4E: [`\u4FB5`].string() // U+4FB5 <cjk>
	0x4F: [`\u5507`].string() // U+5507 <cjk>
	0x50: [`\u5A20`].string() // U+5A20 <cjk>
	0x51: [`\u5BDD`].string() // U+5BDD <cjk>
	0x52: [`\u5BE9`].string() // U+5BE9 <cjk>
	0x53: [`\u5FC3`].string() // U+5FC3 <cjk>
	0x54: [`\u614E`].string() // U+614E <cjk>
	0x55: [`\u632F`].string() // U+632F <cjk>
	0x56: [`\u65B0`].string() // U+65B0 <cjk>
	0x57: [`\u664B`].string() // U+664B <cjk>
	0x58: [`\u68EE`].string() // U+68EE <cjk>
	0x59: [`\u699B`].string() // U+699B <cjk>
	0x5A: [`\u6D78`].string() // U+6D78 <cjk>
	0x5B: [`\u6DF1`].string() // U+6DF1 <cjk>
	0x5C: [`\u7533`].string() // U+7533 <cjk>
	0x5D: [`\u75B9`].string() // U+75B9 <cjk>
	0x5E: [`\u771F`].string() // U+771F <cjk>
	0x5F: [`\u795E`].string() // U+795E <cjk>
	0x60: [`\u79E6`].string() // U+79E6 <cjk>
	0x61: [`\u7D33`].string() // U+7D33 <cjk>
	0x62: [`\u81E3`].string() // U+81E3 <cjk>
	0x63: [`\u82AF`].string() // U+82AF <cjk>
	0x64: [`\u85AA`].string() // U+85AA <cjk>
	0x65: [`\u89AA`].string() // U+89AA <cjk>
	0x66: [`\u8A3A`].string() // U+8A3A <cjk>
	0x67: [`\u8EAB`].string() // U+8EAB <cjk>
	0x68: [`\u8F9B`].string() // U+8F9B <cjk>
	0x69: [`\u9032`].string() // U+9032 <cjk>
	0x6A: [`\u91DD`].string() // U+91DD <cjk>
	0x6B: [`\u9707`].string() // U+9707 <cjk>
	0x6C: [`\u4EBA`].string() // U+4EBA <cjk>
	0x6D: [`\u4EC1`].string() // U+4EC1 <cjk>
	0x6E: [`\u5203`].string() // U+5203 <cjk>
	0x6F: [`\u5875`].string() // U+5875 <cjk>
	0x70: [`\u58EC`].string() // U+58EC <cjk>
	0x71: [`\u5C0B`].string() // U+5C0B <cjk>
	0x72: [`\u751A`].string() // U+751A <cjk>
	0x73: [`\u5C3D`].string() // U+5C3D <cjk>
	0x74: [`\u814E`].string() // U+814E <cjk>
	0x75: [`\u8A0A`].string() // U+8A0A <cjk>
	0x76: [`\u8FC5`].string() // U+8FC5 <cjk>
	0x77: [`\u9663`].string() // U+9663 <cjk>
	0x78: [`\u976D`].string() // U+976D <cjk>
	0x79: [`\u7B25`].string() // U+7B25 <cjk>
	0x7A: [`\u8ACF`].string() // U+8ACF <cjk>
	0x7B: [`\u9808`].string() // U+9808 <cjk>
	0x7C: [`\u9162`].string() // U+9162 <cjk>
	0x7D: [`\u56F3`].string() // U+56F3 <cjk>
	0x7E: [`\u53A8`].string() // U+53A8 <cjk>
	0x80: [`\u9017`].string() // U+9017 <cjk>
	0x81: [`\u5439`].string() // U+5439 <cjk>
	0x82: [`\u5782`].string() // U+5782 <cjk>
	0x83: [`\u5E25`].string() // U+5E25 <cjk>
	0x84: [`\u63A8`].string() // U+63A8 <cjk>
	0x85: [`\u6C34`].string() // U+6C34 <cjk>
	0x86: [`\u708A`].string() // U+708A <cjk>
	0x87: [`\u7761`].string() // U+7761 <cjk>
	0x88: [`\u7C8B`].string() // U+7C8B <cjk>
	0x89: [`\u7FE0`].string() // U+7FE0 <cjk>
	0x8A: [`\u8870`].string() // U+8870 <cjk>
	0x8B: [`\u9042`].string() // U+9042 <cjk>
	0x8C: [`\u9154`].string() // U+9154 <cjk>
	0x8D: [`\u9310`].string() // U+9310 <cjk>
	0x8E: [`\u9318`].string() // U+9318 <cjk>
	0x8F: [`\u968F`].string() // U+968F <cjk>
	0x90: [`\u745E`].string() // U+745E <cjk>
	0x91: [`\u9AC4`].string() // U+9AC4 <cjk>
	0x92: [`\u5D07`].string() // U+5D07 <cjk>
	0x93: [`\u5D69`].string() // U+5D69 <cjk>
	0x94: [`\u6570`].string() // U+6570 <cjk>
	0x95: [`\u67A2`].string() // U+67A2 <cjk>
	0x96: [`\u8DA8`].string() // U+8DA8 <cjk>
	0x97: [`\u96DB`].string() // U+96DB <cjk>
	0x98: [`\u636E`].string() // U+636E <cjk>
	0x99: [`\u6749`].string() // U+6749 <cjk>
	0x9A: [`\u6919`].string() // U+6919 <cjk>
	0x9B: [`\u83C5`].string() // U+83C5 <cjk>
	0x9C: [`\u9817`].string() // U+9817 <cjk>
	0x9D: [`\u96C0`].string() // U+96C0 <cjk>
	0x9E: [`\u88FE`].string() // U+88FE <cjk>
	0x9F: [`\u6F84`].string() // U+6F84 <cjk>
	0xA0: [`\u647A`].string() // U+647A <cjk>
	0xA1: [`\u5BF8`].string() // U+5BF8 <cjk>
	0xA2: [`\u4E16`].string() // U+4E16 <cjk>
	0xA3: [`\u702C`].string() // U+702C <cjk>
	0xA4: [`\u755D`].string() // U+755D <cjk>
	0xA5: [`\u662F`].string() // U+662F <cjk>
	0xA6: [`\u51C4`].string() // U+51C4 <cjk>
	0xA7: [`\u5236`].string() // U+5236 <cjk>
	0xA8: [`\u52E2`].string() // U+52E2 <cjk>
	0xA9: [`\u59D3`].string() // U+59D3 <cjk>
	0xAA: [`\u5F81`].string() // U+5F81 <cjk>
	0xAB: [`\u6027`].string() // U+6027 <cjk>
	0xAC: [`\u6210`].string() // U+6210 <cjk>
	0xAD: [`\u653F`].string() // U+653F <cjk>
	0xAE: [`\u6574`].string() // U+6574 <cjk>
	0xAF: [`\u661F`].string() // U+661F <cjk>
	0xB0: [`\u6674`].string() // U+6674 <cjk>
	0xB1: [`\u68F2`].string() // U+68F2 <cjk>
	0xB2: [`\u6816`].string() // U+6816 <cjk>
	0xB3: [`\u6B63`].string() // U+6B63 <cjk>
	0xB4: [`\u6E05`].string() // U+6E05 <cjk>
	0xB5: [`\u7272`].string() // U+7272 <cjk>
	0xB6: [`\u751F`].string() // U+751F <cjk>
	0xB7: [`\u76DB`].string() // U+76DB <cjk>
	0xB8: [`\u7CBE`].string() // U+7CBE <cjk>
	0xB9: [`\u8056`].string() // U+8056 <cjk>
	0xBA: [`\u58F0`].string() // U+58F0 <cjk>
	0xBB: [`\u88FD`].string() // U+88FD <cjk>
	0xBC: [`\u897F`].string() // U+897F <cjk>
	0xBD: [`\u8AA0`].string() // U+8AA0 <cjk>
	0xBE: [`\u8A93`].string() // U+8A93 <cjk>
	0xBF: [`\u8ACB`].string() // U+8ACB <cjk>
	0xC0: [`\u901D`].string() // U+901D <cjk>
	0xC1: [`\u9192`].string() // U+9192 <cjk>
	0xC2: [`\u9752`].string() // U+9752 <cjk>
	0xC3: [`\u9759`].string() // U+9759 <cjk>
	0xC4: [`\u6589`].string() // U+6589 <cjk>
	0xC5: [`\u7A0E`].string() // U+7A0E <cjk>
	0xC6: [`\u8106`].string() // U+8106 <cjk>
	0xC7: [`\u96BB`].string() // U+96BB <cjk>
	0xC8: [`\u5E2D`].string() // U+5E2D <cjk>
	0xC9: [`\u60DC`].string() // U+60DC <cjk>
	0xCA: [`\u621A`].string() // U+621A <cjk>
	0xCB: [`\u65A5`].string() // U+65A5 <cjk>
	0xCC: [`\u6614`].string() // U+6614 <cjk>
	0xCD: [`\u6790`].string() // U+6790 <cjk>
	0xCE: [`\u77F3`].string() // U+77F3 <cjk>
	0xCF: [`\u7A4D`].string() // U+7A4D <cjk>
	0xD0: [`\u7C4D`].string() // U+7C4D <cjk>
	0xD1: [`\u7E3E`].string() // U+7E3E <cjk>
	0xD2: [`\u810A`].string() // U+810A <cjk>
	0xD3: [`\u8CAC`].string() // U+8CAC <cjk>
	0xD4: [`\u8D64`].string() // U+8D64 <cjk>
	0xD5: [`\u8DE1`].string() // U+8DE1 <cjk>
	0xD6: [`\u8E5F`].string() // U+8E5F <cjk>
	0xD7: [`\u78A9`].string() // U+78A9 <cjk>
	0xD8: [`\u5207`].string() // U+5207 <cjk>
	0xD9: [`\u62D9`].string() // U+62D9 <cjk>
	0xDA: [`\u63A5`].string() // U+63A5 <cjk>
	0xDB: [`\u6442`].string() // U+6442 <cjk>
	0xDC: [`\u6298`].string() // U+6298 <cjk>
	0xDD: [`\u8A2D`].string() // U+8A2D <cjk>
	0xDE: [`\u7A83`].string() // U+7A83 <cjk>
	0xDF: [`\u7BC0`].string() // U+7BC0 <cjk>
	0xE0: [`\u8AAC`].string() // U+8AAC <cjk>
	0xE1: [`\u96EA`].string() // U+96EA <cjk>
	0xE2: [`\u7D76`].string() // U+7D76 <cjk>
	0xE3: [`\u820C`].string() // U+820C <cjk>
	0xE4: [`\u8749`].string() // U+8749 <cjk>
	0xE5: [`\u4ED9`].string() // U+4ED9 <cjk>
	0xE6: [`\u5148`].string() // U+5148 <cjk>
	0xE7: [`\u5343`].string() // U+5343 <cjk>
	0xE8: [`\u5360`].string() // U+5360 <cjk>
	0xE9: [`\u5BA3`].string() // U+5BA3 <cjk>
	0xEA: [`\u5C02`].string() // U+5C02 <cjk>
	0xEB: [`\u5C16`].string() // U+5C16 <cjk>
	0xEC: [`\u5DDD`].string() // U+5DDD <cjk>
	0xED: [`\u6226`].string() // U+6226 <cjk>
	0xEE: [`\u6247`].string() // U+6247 <cjk>
	0xEF: [`\u64B0`].string() // U+64B0 <cjk>
	0xF0: [`\u6813`].string() // U+6813 <cjk>
	0xF1: [`\u6834`].string() // U+6834 <cjk>
	0xF2: [`\u6CC9`].string() // U+6CC9 <cjk>
	0xF3: [`\u6D45`].string() // U+6D45 <cjk>
	0xF4: [`\u6D17`].string() // U+6D17 <cjk>
	0xF5: [`\u67D3`].string() // U+67D3 <cjk>
	0xF6: [`\u6F5C`].string() // U+6F5C <cjk>
	0xF7: [`\u714E`].string() // U+714E <cjk>
	0xF8: [`\u717D`].string() // U+717D <cjk>
	0xF9: [`\u65CB`].string() // U+65CB <cjk>
	0xFA: [`\u7A7F`].string() // U+7A7F <cjk>
	0xFB: [`\u7BAD`].string() // U+7BAD <cjk>
	0xFC: [`\u7DDA`].string() // U+7DDA <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x87 = {
	0x40: [`\u2460`].string() // U+2460 CIRCLED DIGIT ONE
	0x41: [`\u2461`].string() // U+2461 CIRCLED DIGIT TWO
	0x42: [`\u2462`].string() // U+2462 CIRCLED DIGIT THREE
	0x43: [`\u2463`].string() // U+2463 CIRCLED DIGIT FOUR
	0x44: [`\u2464`].string() // U+2464 CIRCLED DIGIT FIVE
	0x45: [`\u2465`].string() // U+2465 CIRCLED DIGIT SIX
	0x46: [`\u2466`].string() // U+2466 CIRCLED DIGIT SEVEN
	0x47: [`\u2467`].string() // U+2467 CIRCLED DIGIT EIGHT
	0x48: [`\u2468`].string() // U+2468 CIRCLED DIGIT NINE
	0x49: [`\u2469`].string() // U+2469 CIRCLED NUMBER TEN
	0x4A: [`\u246A`].string() // U+246A CIRCLED NUMBER ELEVEN
	0x4B: [`\u246B`].string() // U+246B CIRCLED NUMBER TWELVE
	0x4C: [`\u246C`].string() // U+246C CIRCLED NUMBER THIRTEEN
	0x4D: [`\u246D`].string() // U+246D CIRCLED NUMBER FOURTEEN
	0x4E: [`\u246E`].string() // U+246E CIRCLED NUMBER FIFTEEN
	0x4F: [`\u246F`].string() // U+246F CIRCLED NUMBER SIXTEEN
	0x50: [`\u2470`].string() // U+2470 CIRCLED NUMBER SEVENTEEN
	0x51: [`\u2471`].string() // U+2471 CIRCLED NUMBER EIGHTEEN
	0x52: [`\u2472`].string() // U+2472 CIRCLED NUMBER NINETEEN
	0x53: [`\u2473`].string() // U+2473 CIRCLED NUMBER TWENTY
	0x54: [`\u2160`].string() // U+2160 ROMAN NUMERAL ONE
	0x55: [`\u2161`].string() // U+2161 ROMAN NUMERAL TWO
	0x56: [`\u2162`].string() // U+2162 ROMAN NUMERAL THREE
	0x57: [`\u2163`].string() // U+2163 ROMAN NUMERAL FOUR
	0x58: [`\u2164`].string() // U+2164 ROMAN NUMERAL FIVE
	0x59: [`\u2165`].string() // U+2165 ROMAN NUMERAL SIX
	0x5A: [`\u2166`].string() // U+2166 ROMAN NUMERAL SEVEN
	0x5B: [`\u2167`].string() // U+2167 ROMAN NUMERAL EIGHT
	0x5C: [`\u2168`].string() // U+2168 ROMAN NUMERAL NINE
	0x5D: [`\u2169`].string() // U+2169 ROMAN NUMERAL TEN
	0x5E: [`\u216A`].string() // U+216A ROMAN NUMERAL ELEVEN
	0x5F: [`\u3349`].string() // U+3349 SQUARE MIRI
	0x60: [`\u3314`].string() // U+3314 SQUARE KIRO
	0x61: [`\u3322`].string() // U+3322 SQUARE SENTI
	0x62: [`\u334D`].string() // U+334D SQUARE MEETORU
	0x63: [`\u3318`].string() // U+3318 SQUARE GURAMU
	0x64: [`\u3327`].string() // U+3327 SQUARE TON
	0x65: [`\u3303`].string() // U+3303 SQUARE AARU
	0x66: [`\u3336`].string() // U+3336 SQUARE HEKUTAARU
	0x67: [`\u3351`].string() // U+3351 SQUARE RITTORU
	0x68: [`\u3357`].string() // U+3357 SQUARE WATTO
	0x69: [`\u330D`].string() // U+330D SQUARE KARORII
	0x6A: [`\u3326`].string() // U+3326 SQUARE DORU
	0x6B: [`\u3323`].string() // U+3323 SQUARE SENTO
	0x6C: [`\u332B`].string() // U+332B SQUARE PAASENTO
	0x6D: [`\u334A`].string() // U+334A SQUARE MIRIBAARU
	0x6E: [`\u333B`].string() // U+333B SQUARE PEEZI
	0x6F: [`\u339C`].string() // U+339C SQUARE MM
	0x70: [`\u339D`].string() // U+339D SQUARE CM
	0x71: [`\u339E`].string() // U+339E SQUARE KM
	0x72: [`\u338E`].string() // U+338E SQUARE MG
	0x73: [`\u338F`].string() // U+338F SQUARE KG
	0x74: [`\u33C4`].string() // U+33C4 SQUARE CC
	0x75: [`\u33A1`].string() // U+33A1 SQUARE M SQUARED
	0x76: [`\u216B`].string() // U+216B ROMAN NUMERAL TWELVE
	0x7E: [`\u337B`].string() // U+337B SQUARE ERA NAME HEISEI
	0x80: [`\u301D`].string() // U+301D REVERSED DOUBLE PRIME QUOTATION MARK
	0x81: [`\u301F`].string() // U+301F LOW DOUBLE PRIME QUOTATION MARK
	0x82: [`\u2116`].string() // U+2116 NUMERO SIGN
	0x83: [`\u33CD`].string() // U+33CD SQUARE KK
	0x84: [`\u2121`].string() // U+2121 TELEPHONE SIGN
	0x85: [`\u32A4`].string() // U+32A4 CIRCLED IDEOGRAPH HIGH
	0x86: [`\u32A5`].string() // U+32A5 CIRCLED IDEOGRAPH CENTRE
	0x87: [`\u32A6`].string() // U+32A6 CIRCLED IDEOGRAPH LOW
	0x88: [`\u32A7`].string() // U+32A7 CIRCLED IDEOGRAPH LEFT
	0x89: [`\u32A8`].string() // U+32A8 CIRCLED IDEOGRAPH RIGHT
	0x8A: [`\u3231`].string() // U+3231 PARENTHESIZED IDEOGRAPH STOCK
	0x8B: [`\u3232`].string() // U+3232 PARENTHESIZED IDEOGRAPH HAVE
	0x8C: [`\u3239`].string() // U+3239 PARENTHESIZED IDEOGRAPH REPRESENT
	0x8D: [`\u337E`].string() // U+337E SQUARE ERA NAME MEIZI
	0x8E: [`\u337D`].string() // U+337D SQUARE ERA NAME TAISYOU
	0x8F: [`\u337C`].string() // U+337C SQUARE ERA NAME SYOUWA
	0x93: [`\u222E`].string() // U+222E CONTOUR INTEGRAL
	0x98: [`\u221F`].string() // U+221F RIGHT ANGLE
	0x99: [`\u22BF`].string() // U+22BF RIGHT TRIANGLE
	0x9D: [`\u2756`].string() // U+2756 BLACK DIAMOND MINUS WHITE X
	0x9E: [`\u261E`].string() // U+261E WHITE RIGHT POINTING INDEX
	0x9F: [`\u4FF1`].string() // U+4FF1 <cjk>
	0xA0: utf32_to_str(0x2000B) // U+2000B <cjk>
	0xA1: [`\u3402`].string() // U+3402 <cjk>
	0xA2: [`\u4E28`].string() // U+4E28 <cjk>
	0xA3: [`\u4E2F`].string() // U+4E2F <cjk>
	0xA4: [`\u4E30`].string() // U+4E30 <cjk>
	0xA5: [`\u4E8D`].string() // U+4E8D <cjk>
	0xA6: [`\u4EE1`].string() // U+4EE1 <cjk>
	0xA7: [`\u4EFD`].string() // U+4EFD <cjk>
	0xA8: [`\u4EFF`].string() // U+4EFF <cjk>
	0xA9: [`\u4F03`].string() // U+4F03 <cjk>
	0xAA: [`\u4F0B`].string() // U+4F0B <cjk>
	0xAB: [`\u4F60`].string() // U+4F60 <cjk>
	0xAC: [`\u4F48`].string() // U+4F48 <cjk>
	0xAD: [`\u4F49`].string() // U+4F49 <cjk>
	0xAE: [`\u4F56`].string() // U+4F56 <cjk>
	0xAF: [`\u4F5F`].string() // U+4F5F <cjk>
	0xB0: [`\u4F6A`].string() // U+4F6A <cjk>
	0xB1: [`\u4F6C`].string() // U+4F6C <cjk>
	0xB2: [`\u4F7E`].string() // U+4F7E <cjk>
	0xB3: [`\u4F8A`].string() // U+4F8A <cjk>
	0xB4: [`\u4F94`].string() // U+4F94 <cjk>
	0xB5: [`\u4F97`].string() // U+4F97 <cjk>
	0xB6: [`\uFA30`].string() // U+FA30 CJK COMPATIBILITY IDEOGRAPH-FA30
	0xB7: [`\u4FC9`].string() // U+4FC9 <cjk>
	0xB8: [`\u4FE0`].string() // U+4FE0 <cjk>
	0xB9: [`\u5001`].string() // U+5001 <cjk>
	0xBA: [`\u5002`].string() // U+5002 <cjk>
	0xBB: [`\u500E`].string() // U+500E <cjk>
	0xBC: [`\u5018`].string() // U+5018 <cjk>
	0xBD: [`\u5027`].string() // U+5027 <cjk>
	0xBE: [`\u502E`].string() // U+502E <cjk>
	0xBF: [`\u5040`].string() // U+5040 <cjk>
	0xC0: [`\u503B`].string() // U+503B <cjk>
	0xC1: [`\u5041`].string() // U+5041 <cjk>
	0xC2: [`\u5094`].string() // U+5094 <cjk>
	0xC3: [`\u50CC`].string() // U+50CC <cjk>
	0xC4: [`\u50F2`].string() // U+50F2 <cjk>
	0xC5: [`\u50D0`].string() // U+50D0 <cjk>
	0xC6: [`\u50E6`].string() // U+50E6 <cjk>
	0xC7: [`\uFA31`].string() // U+FA31 CJK COMPATIBILITY IDEOGRAPH-FA31
	0xC8: [`\u5106`].string() // U+5106 <cjk>
	0xC9: [`\u5103`].string() // U+5103 <cjk>
	0xCA: [`\u510B`].string() // U+510B <cjk>
	0xCB: [`\u511E`].string() // U+511E <cjk>
	0xCC: [`\u5135`].string() // U+5135 <cjk>
	0xCD: [`\u514A`].string() // U+514A <cjk>
	0xCE: [`\uFA32`].string() // U+FA32 CJK COMPATIBILITY IDEOGRAPH-FA32
	0xCF: [`\u5155`].string() // U+5155 <cjk>
	0xD0: [`\u5157`].string() // U+5157 <cjk>
	0xD1: [`\u34B5`].string() // U+34B5 <cjk>
	0xD2: [`\u519D`].string() // U+519D <cjk>
	0xD3: [`\u51C3`].string() // U+51C3 <cjk>
	0xD4: [`\u51CA`].string() // U+51CA <cjk>
	0xD5: [`\u51DE`].string() // U+51DE <cjk>
	0xD6: [`\u51E2`].string() // U+51E2 <cjk>
	0xD7: [`\u51EE`].string() // U+51EE <cjk>
	0xD8: [`\u5201`].string() // U+5201 <cjk>
	0xD9: [`\u34DB`].string() // U+34DB <cjk>
	0xDA: [`\u5213`].string() // U+5213 <cjk>
	0xDB: [`\u5215`].string() // U+5215 <cjk>
	0xDC: [`\u5249`].string() // U+5249 <cjk>
	0xDD: [`\u5257`].string() // U+5257 <cjk>
	0xDE: [`\u5261`].string() // U+5261 <cjk>
	0xDF: [`\u5293`].string() // U+5293 <cjk>
	0xE0: [`\u52C8`].string() // U+52C8 <cjk>
	0xE1: [`\uFA33`].string() // U+FA33 CJK COMPATIBILITY IDEOGRAPH-FA33
	0xE2: [`\u52CC`].string() // U+52CC <cjk>
	0xE3: [`\u52D0`].string() // U+52D0 <cjk>
	0xE4: [`\u52D6`].string() // U+52D6 <cjk>
	0xE5: [`\u52DB`].string() // U+52DB <cjk>
	0xE6: [`\uFA34`].string() // U+FA34 CJK COMPATIBILITY IDEOGRAPH-FA34
	0xE7: [`\u52F0`].string() // U+52F0 <cjk>
	0xE8: [`\u52FB`].string() // U+52FB <cjk>
	0xE9: [`\u5300`].string() // U+5300 <cjk>
	0xEA: [`\u5307`].string() // U+5307 <cjk>
	0xEB: [`\u531C`].string() // U+531C <cjk>
	0xEC: [`\uFA35`].string() // U+FA35 CJK COMPATIBILITY IDEOGRAPH-FA35
	0xED: [`\u5361`].string() // U+5361 <cjk>
	0xEE: [`\u5363`].string() // U+5363 <cjk>
	0xEF: [`\u537D`].string() // U+537D <cjk>
	0xF0: [`\u5393`].string() // U+5393 <cjk>
	0xF1: [`\u539D`].string() // U+539D <cjk>
	0xF2: [`\u53B2`].string() // U+53B2 <cjk>
	0xF3: [`\u5412`].string() // U+5412 <cjk>
	0xF4: [`\u5427`].string() // U+5427 <cjk>
	0xF5: [`\u544D`].string() // U+544D <cjk>
	0xF6: [`\u549C`].string() // U+549C <cjk>
	0xF7: [`\u546B`].string() // U+546B <cjk>
	0xF8: [`\u5474`].string() // U+5474 <cjk>
	0xF9: [`\u547F`].string() // U+547F <cjk>
	0xFA: [`\u5488`].string() // U+5488 <cjk>
	0xFB: [`\u5496`].string() // U+5496 <cjk>
	0xFC: [`\u54A1`].string() // U+54A1 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x93 = {
	0x40: [`\u90B8`].string() // U+90B8 <cjk>
	0x41: [`\u912D`].string() // U+912D <cjk>
	0x42: [`\u91D8`].string() // U+91D8 <cjk>
	0x43: [`\u9F0E`].string() // U+9F0E <cjk>
	0x44: [`\u6CE5`].string() // U+6CE5 <cjk>
	0x45: [`\u6458`].string() // U+6458 <cjk>
	0x46: [`\u64E2`].string() // U+64E2 <cjk>
	0x47: [`\u6575`].string() // U+6575 <cjk>
	0x48: [`\u6EF4`].string() // U+6EF4 <cjk>
	0x49: [`\u7684`].string() // U+7684 <cjk>
	0x4A: [`\u7B1B`].string() // U+7B1B <cjk>
	0x4B: [`\u9069`].string() // U+9069 <cjk>
	0x4C: [`\u93D1`].string() // U+93D1 <cjk>
	0x4D: [`\u6EBA`].string() // U+6EBA <cjk>
	0x4E: [`\u54F2`].string() // U+54F2 <cjk>
	0x4F: [`\u5FB9`].string() // U+5FB9 <cjk>
	0x50: [`\u64A4`].string() // U+64A4 <cjk>
	0x51: [`\u8F4D`].string() // U+8F4D <cjk>
	0x52: [`\u8FED`].string() // U+8FED <cjk>
	0x53: [`\u9244`].string() // U+9244 <cjk>
	0x54: [`\u5178`].string() // U+5178 <cjk>
	0x55: [`\u586B`].string() // U+586B <cjk>
	0x56: [`\u5929`].string() // U+5929 <cjk>
	0x57: [`\u5C55`].string() // U+5C55 <cjk>
	0x58: [`\u5E97`].string() // U+5E97 <cjk>
	0x59: [`\u6DFB`].string() // U+6DFB <cjk>
	0x5A: [`\u7E8F`].string() // U+7E8F <cjk>
	0x5B: [`\u751C`].string() // U+751C <cjk>
	0x5C: [`\u8CBC`].string() // U+8CBC <cjk>
	0x5D: [`\u8EE2`].string() // U+8EE2 <cjk>
	0x5E: [`\u985B`].string() // U+985B <cjk>
	0x5F: [`\u70B9`].string() // U+70B9 <cjk>
	0x60: [`\u4F1D`].string() // U+4F1D <cjk>
	0x61: [`\u6BBF`].string() // U+6BBF <cjk>
	0x62: [`\u6FB1`].string() // U+6FB1 <cjk>
	0x63: [`\u7530`].string() // U+7530 <cjk>
	0x64: [`\u96FB`].string() // U+96FB <cjk>
	0x65: [`\u514E`].string() // U+514E <cjk>
	0x66: [`\u5410`].string() // U+5410 <cjk>
	0x67: [`\u5835`].string() // U+5835 <cjk>
	0x68: [`\u5857`].string() // U+5857 <cjk>
	0x69: [`\u59AC`].string() // U+59AC <cjk>
	0x6A: [`\u5C60`].string() // U+5C60 <cjk>
	0x6B: [`\u5F92`].string() // U+5F92 <cjk>
	0x6C: [`\u6597`].string() // U+6597 <cjk>
	0x6D: [`\u675C`].string() // U+675C <cjk>
	0x6E: [`\u6E21`].string() // U+6E21 <cjk>
	0x6F: [`\u767B`].string() // U+767B <cjk>
	0x70: [`\u83DF`].string() // U+83DF <cjk>
	0x71: [`\u8CED`].string() // U+8CED <cjk>
	0x72: [`\u9014`].string() // U+9014 <cjk>
	0x73: [`\u90FD`].string() // U+90FD <cjk>
	0x74: [`\u934D`].string() // U+934D <cjk>
	0x75: [`\u7825`].string() // U+7825 <cjk>
	0x76: [`\u783A`].string() // U+783A <cjk>
	0x77: [`\u52AA`].string() // U+52AA <cjk>
	0x78: [`\u5EA6`].string() // U+5EA6 <cjk>
	0x79: [`\u571F`].string() // U+571F <cjk>
	0x7A: [`\u5974`].string() // U+5974 <cjk>
	0x7B: [`\u6012`].string() // U+6012 <cjk>
	0x7C: [`\u5012`].string() // U+5012 <cjk>
	0x7D: [`\u515A`].string() // U+515A <cjk>
	0x7E: [`\u51AC`].string() // U+51AC <cjk>
	0x80: [`\u51CD`].string() // U+51CD <cjk>
	0x81: [`\u5200`].string() // U+5200 <cjk>
	0x82: [`\u5510`].string() // U+5510 <cjk>
	0x83: [`\u5854`].string() // U+5854 <cjk>
	0x84: [`\u5858`].string() // U+5858 <cjk>
	0x85: [`\u5957`].string() // U+5957 <cjk>
	0x86: [`\u5B95`].string() // U+5B95 <cjk>
	0x87: [`\u5CF6`].string() // U+5CF6 <cjk>
	0x88: [`\u5D8B`].string() // U+5D8B <cjk>
	0x89: [`\u60BC`].string() // U+60BC <cjk>
	0x8A: [`\u6295`].string() // U+6295 <cjk>
	0x8B: [`\u642D`].string() // U+642D <cjk>
	0x8C: [`\u6771`].string() // U+6771 <cjk>
	0x8D: [`\u6843`].string() // U+6843 <cjk>
	0x8E: [`\u68BC`].string() // U+68BC <cjk>
	0x8F: [`\u68DF`].string() // U+68DF <cjk>
	0x90: [`\u76D7`].string() // U+76D7 <cjk>
	0x91: [`\u6DD8`].string() // U+6DD8 <cjk>
	0x92: [`\u6E6F`].string() // U+6E6F <cjk>
	0x93: [`\u6D9B`].string() // U+6D9B <cjk>
	0x94: [`\u706F`].string() // U+706F <cjk>
	0x95: [`\u71C8`].string() // U+71C8 <cjk>
	0x96: [`\u5F53`].string() // U+5F53 <cjk>
	0x97: [`\u75D8`].string() // U+75D8 <cjk>
	0x98: [`\u7977`].string() // U+7977 <cjk>
	0x99: [`\u7B49`].string() // U+7B49 <cjk>
	0x9A: [`\u7B54`].string() // U+7B54 <cjk>
	0x9B: [`\u7B52`].string() // U+7B52 <cjk>
	0x9C: [`\u7CD6`].string() // U+7CD6 <cjk>
	0x9D: [`\u7D71`].string() // U+7D71 <cjk>
	0x9E: [`\u5230`].string() // U+5230 <cjk>
	0x9F: [`\u8463`].string() // U+8463 <cjk>
	0xA0: [`\u8569`].string() // U+8569 <cjk>
	0xA1: [`\u85E4`].string() // U+85E4 <cjk>
	0xA2: [`\u8A0E`].string() // U+8A0E <cjk>
	0xA3: [`\u8B04`].string() // U+8B04 <cjk>
	0xA4: [`\u8C46`].string() // U+8C46 <cjk>
	0xA5: [`\u8E0F`].string() // U+8E0F <cjk>
	0xA6: [`\u9003`].string() // U+9003 <cjk>
	0xA7: [`\u900F`].string() // U+900F <cjk>
	0xA8: [`\u9419`].string() // U+9419 <cjk>
	0xA9: [`\u9676`].string() // U+9676 <cjk>
	0xAA: [`\u982D`].string() // U+982D <cjk>
	0xAB: [`\u9A30`].string() // U+9A30 <cjk>
	0xAC: [`\u95D8`].string() // U+95D8 <cjk>
	0xAD: [`\u50CD`].string() // U+50CD <cjk>
	0xAE: [`\u52D5`].string() // U+52D5 <cjk>
	0xAF: [`\u540C`].string() // U+540C <cjk>
	0xB0: [`\u5802`].string() // U+5802 <cjk>
	0xB1: [`\u5C0E`].string() // U+5C0E <cjk>
	0xB2: [`\u61A7`].string() // U+61A7 <cjk>
	0xB3: [`\u649E`].string() // U+649E <cjk>
	0xB4: [`\u6D1E`].string() // U+6D1E <cjk>
	0xB5: [`\u77B3`].string() // U+77B3 <cjk>
	0xB6: [`\u7AE5`].string() // U+7AE5 <cjk>
	0xB7: [`\u80F4`].string() // U+80F4 <cjk>
	0xB8: [`\u8404`].string() // U+8404 <cjk>
	0xB9: [`\u9053`].string() // U+9053 <cjk>
	0xBA: [`\u9285`].string() // U+9285 <cjk>
	0xBB: [`\u5CE0`].string() // U+5CE0 <cjk>
	0xBC: [`\u9D07`].string() // U+9D07 <cjk>
	0xBD: [`\u533F`].string() // U+533F <cjk>
	0xBE: [`\u5F97`].string() // U+5F97 <cjk>
	0xBF: [`\u5FB3`].string() // U+5FB3 <cjk>
	0xC0: [`\u6D9C`].string() // U+6D9C <cjk>
	0xC1: [`\u7279`].string() // U+7279 <cjk>
	0xC2: [`\u7763`].string() // U+7763 <cjk>
	0xC3: [`\u79BF`].string() // U+79BF <cjk>
	0xC4: [`\u7BE4`].string() // U+7BE4 <cjk>
	0xC5: [`\u6BD2`].string() // U+6BD2 <cjk>
	0xC6: [`\u72EC`].string() // U+72EC <cjk>
	0xC7: [`\u8AAD`].string() // U+8AAD <cjk>
	0xC8: [`\u6803`].string() // U+6803 <cjk>
	0xC9: [`\u6A61`].string() // U+6A61 <cjk>
	0xCA: [`\u51F8`].string() // U+51F8 <cjk>
	0xCB: [`\u7A81`].string() // U+7A81 <cjk>
	0xCC: [`\u6934`].string() // U+6934 <cjk>
	0xCD: [`\u5C4A`].string() // U+5C4A <cjk>
	0xCE: [`\u9CF6`].string() // U+9CF6 <cjk>
	0xCF: [`\u82EB`].string() // U+82EB <cjk>
	0xD0: [`\u5BC5`].string() // U+5BC5 <cjk>
	0xD1: [`\u9149`].string() // U+9149 <cjk>
	0xD2: [`\u701E`].string() // U+701E <cjk>
	0xD3: [`\u5678`].string() // U+5678 <cjk>
	0xD4: [`\u5C6F`].string() // U+5C6F <cjk>
	0xD5: [`\u60C7`].string() // U+60C7 <cjk>
	0xD6: [`\u6566`].string() // U+6566 <cjk>
	0xD7: [`\u6C8C`].string() // U+6C8C <cjk>
	0xD8: [`\u8C5A`].string() // U+8C5A <cjk>
	0xD9: [`\u9041`].string() // U+9041 <cjk>
	0xDA: [`\u9813`].string() // U+9813 <cjk>
	0xDB: [`\u5451`].string() // U+5451 <cjk>
	0xDC: [`\u66C7`].string() // U+66C7 <cjk>
	0xDD: [`\u920D`].string() // U+920D <cjk>
	0xDE: [`\u5948`].string() // U+5948 <cjk>
	0xDF: [`\u90A3`].string() // U+90A3 <cjk>
	0xE0: [`\u5185`].string() // U+5185 <cjk>
	0xE1: [`\u4E4D`].string() // U+4E4D <cjk>
	0xE2: [`\u51EA`].string() // U+51EA <cjk>
	0xE3: [`\u8599`].string() // U+8599 <cjk>
	0xE4: [`\u8B0E`].string() // U+8B0E <cjk>
	0xE5: [`\u7058`].string() // U+7058 <cjk>
	0xE6: [`\u637A`].string() // U+637A <cjk>
	0xE7: [`\u934B`].string() // U+934B <cjk>
	0xE8: [`\u6962`].string() // U+6962 <cjk>
	0xE9: [`\u99B4`].string() // U+99B4 <cjk>
	0xEA: [`\u7E04`].string() // U+7E04 <cjk>
	0xEB: [`\u7577`].string() // U+7577 <cjk>
	0xEC: [`\u5357`].string() // U+5357 <cjk>
	0xED: [`\u6960`].string() // U+6960 <cjk>
	0xEE: [`\u8EDF`].string() // U+8EDF <cjk>
	0xEF: [`\u96E3`].string() // U+96E3 <cjk>
	0xF0: [`\u6C5D`].string() // U+6C5D <cjk>
	0xF1: [`\u4E8C`].string() // U+4E8C <cjk>
	0xF2: [`\u5C3C`].string() // U+5C3C <cjk>
	0xF3: [`\u5F10`].string() // U+5F10 <cjk>
	0xF4: [`\u8FE9`].string() // U+8FE9 <cjk>
	0xF5: [`\u5302`].string() // U+5302 <cjk>
	0xF6: [`\u8CD1`].string() // U+8CD1 <cjk>
	0xF7: [`\u8089`].string() // U+8089 <cjk>
	0xF8: [`\u8679`].string() // U+8679 <cjk>
	0xF9: [`\u5EFF`].string() // U+5EFF <cjk>
	0xFA: [`\u65E5`].string() // U+65E5 <cjk>
	0xFB: [`\u4E73`].string() // U+4E73 <cjk>
	0xFC: [`\u5165`].string() // U+5165 <cjk>
}

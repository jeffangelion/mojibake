module mojibake

const utf8_to_jis_x_0213_data = {
	`¥`: [u8(0x5C)] // U+00A5 YEN SIGN
	`‾`: [u8(0x7E)] // U+203E OVERLINE
	`｡`: [u8(0xA1)] // U+FF61 HALFWIDTH IDEOGRAPHIC FULL STOP
	`｢`: [u8(0xA2)] // U+FF62 HALFWIDTH LEFT CORNER BRACKET
	`｣`: [u8(0xA3)] // U+FF63 HALFWIDTH RIGHT CORNER BRACKET
	`､`: [u8(0xA4)] // U+FF64 HALFWIDTH IDEOGRAPHIC COMMA
	`･`: [u8(0xA5)] // U+FF65 HALFWIDTH KATAKANA MIDDLE DOT
	`ｦ`: [u8(0xA6)] // U+FF66 HALFWIDTH KATAKANA LETTER WO
	`ｧ`: [u8(0xA7)] // U+FF67 HALFWIDTH KATAKANA LETTER SMALL A
	`ｨ`: [u8(0xA8)] // U+FF68 HALFWIDTH KATAKANA LETTER SMALL I
	`ｩ`: [u8(0xA9)] // U+FF69 HALFWIDTH KATAKANA LETTER SMALL U
	`ｪ`: [u8(0xAA)] // U+FF6A HALFWIDTH KATAKANA LETTER SMALL E
	`ｫ`: [u8(0xAB)] // U+FF6B HALFWIDTH KATAKANA LETTER SMALL O
	`ｬ`: [u8(0xAC)] // U+FF6C HALFWIDTH KATAKANA LETTER SMALL YA
	`ｭ`: [u8(0xAD)] // U+FF6D HALFWIDTH KATAKANA LETTER SMALL YU
	`ｮ`: [u8(0xAE)] // U+FF6E HALFWIDTH KATAKANA LETTER SMALL YO
	`ｯ`: [u8(0xAF)] // U+FF6F HALFWIDTH KATAKANA LETTER SMALL TU
	`ｰ`: [u8(0xB0)] // U+FF70 HALFWIDTH KATAKANA-HIRAGANA PROLONGED SOUND MARK
	`ｱ`: [u8(0xB1)] // U+FF71 HALFWIDTH KATAKANA LETTER A
	`ｲ`: [u8(0xB2)] // U+FF72 HALFWIDTH KATAKANA LETTER I
	`ｳ`: [u8(0xB3)] // U+FF73 HALFWIDTH KATAKANA LETTER U
	`ｴ`: [u8(0xB4)] // U+FF74 HALFWIDTH KATAKANA LETTER E
	`ｵ`: [u8(0xB5)] // U+FF75 HALFWIDTH KATAKANA LETTER O
	`ｶ`: [u8(0xB6)] // U+FF76 HALFWIDTH KATAKANA LETTER KA
	`ｷ`: [u8(0xB7)] // U+FF77 HALFWIDTH KATAKANA LETTER KI
	`ｸ`: [u8(0xB8)] // U+FF78 HALFWIDTH KATAKANA LETTER KU
	`ｹ`: [u8(0xB9)] // U+FF79 HALFWIDTH KATAKANA LETTER KE
	`ｺ`: [u8(0xBA)] // U+FF7A HALFWIDTH KATAKANA LETTER KO
	`ｻ`: [u8(0xBB)] // U+FF7B HALFWIDTH KATAKANA LETTER SA
	`ｼ`: [u8(0xBC)] // U+FF7C HALFWIDTH KATAKANA LETTER SI
	`ｽ`: [u8(0xBD)] // U+FF7D HALFWIDTH KATAKANA LETTER SU
	`ｾ`: [u8(0xBE)] // U+FF7E HALFWIDTH KATAKANA LETTER SE
	`ｿ`: [u8(0xBF)] // U+FF7F HALFWIDTH KATAKANA LETTER SO
	`ﾀ`: [u8(0xC0)] // U+FF80 HALFWIDTH KATAKANA LETTER TA
	`ﾁ`: [u8(0xC1)] // U+FF81 HALFWIDTH KATAKANA LETTER TI
	`ﾂ`: [u8(0xC2)] // U+FF82 HALFWIDTH KATAKANA LETTER TU
	`ﾃ`: [u8(0xC3)] // U+FF83 HALFWIDTH KATAKANA LETTER TE
	`ﾄ`: [u8(0xC4)] // U+FF84 HALFWIDTH KATAKANA LETTER TO
	`ﾅ`: [u8(0xC5)] // U+FF85 HALFWIDTH KATAKANA LETTER NA
	`ﾆ`: [u8(0xC6)] // U+FF86 HALFWIDTH KATAKANA LETTER NI
	`ﾇ`: [u8(0xC7)] // U+FF87 HALFWIDTH KATAKANA LETTER NU
	`ﾈ`: [u8(0xC8)] // U+FF88 HALFWIDTH KATAKANA LETTER NE
	`ﾉ`: [u8(0xC9)] // U+FF89 HALFWIDTH KATAKANA LETTER NO
	`ﾊ`: [u8(0xCA)] // U+FF8A HALFWIDTH KATAKANA LETTER HA
	`ﾋ`: [u8(0xCB)] // U+FF8B HALFWIDTH KATAKANA LETTER HI
	`ﾌ`: [u8(0xCC)] // U+FF8C HALFWIDTH KATAKANA LETTER HU
	`ﾍ`: [u8(0xCD)] // U+FF8D HALFWIDTH KATAKANA LETTER HE
	`ﾎ`: [u8(0xCE)] // U+FF8E HALFWIDTH KATAKANA LETTER HO
	`ﾏ`: [u8(0xCF)] // U+FF8F HALFWIDTH KATAKANA LETTER MA
	`ﾐ`: [u8(0xD0)] // U+FF90 HALFWIDTH KATAKANA LETTER MI
	`ﾑ`: [u8(0xD1)] // U+FF91 HALFWIDTH KATAKANA LETTER MU
	`ﾒ`: [u8(0xD2)] // U+FF92 HALFWIDTH KATAKANA LETTER ME
	`ﾓ`: [u8(0xD3)] // U+FF93 HALFWIDTH KATAKANA LETTER MO
	`ﾔ`: [u8(0xD4)] // U+FF94 HALFWIDTH KATAKANA LETTER YA
	`ﾕ`: [u8(0xD5)] // U+FF95 HALFWIDTH KATAKANA LETTER YU
	`ﾖ`: [u8(0xD6)] // U+FF96 HALFWIDTH KATAKANA LETTER YO
	`ﾗ`: [u8(0xD7)] // U+FF97 HALFWIDTH KATAKANA LETTER RA
	`ﾘ`: [u8(0xD8)] // U+FF98 HALFWIDTH KATAKANA LETTER RI
	`ﾙ`: [u8(0xD9)] // U+FF99 HALFWIDTH KATAKANA LETTER RU
	`ﾚ`: [u8(0xDA)] // U+FF9A HALFWIDTH KATAKANA LETTER RE
	`ﾛ`: [u8(0xDB)] // U+FF9B HALFWIDTH KATAKANA LETTER RO
	`ﾜ`: [u8(0xDC)] // U+FF9C HALFWIDTH KATAKANA LETTER WA
	`ﾝ`: [u8(0xDD)] // U+FF9D HALFWIDTH KATAKANA LETTER N
	`ﾞ`: [u8(0xDE)] // U+FF9E HALFWIDTH KATAKANA VOICED SOUND MARK
	`ﾟ`: [u8(0xDF)] // U+FF9F HALFWIDTH KATAKANA SEMI-VOICED SOUND MARK
	`　`: [u8(0x81), 0x40] // U+3000 IDEOGRAPHIC SPACE
	`、`: [u8(0x81), 0x41] // U+3001 IDEOGRAPHIC COMMA
	`。`: [u8(0x81), 0x42] // U+3002 IDEOGRAPHIC FULL STOP
	`，`: [u8(0x81), 0x43] // U+FF0C FULLWIDTH COMMA
	`．`: [u8(0x81), 0x44] // U+FF0E FULLWIDTH FULL STOP
	`・`: [u8(0x81), 0x45] // U+30FB KATAKANA MIDDLE DOT
	`：`: [u8(0x81), 0x46] // U+FF1A FULLWIDTH COLON
	`；`: [u8(0x81), 0x47] // U+FF1B FULLWIDTH SEMICOLON
	`？`: [u8(0x81), 0x48] // U+FF1F FULLWIDTH QUESTION MARK
	`！`: [u8(0x81), 0x49] // U+FF01 FULLWIDTH EXCLAMATION MARK
	`゛`: [u8(0x81), 0x4A] // U+309B KATAKANA-HIRAGANA VOICED SOUND MARK
	`゜`: [u8(0x81), 0x4B] // U+309C KATAKANA-HIRAGANA SEMI-VOICED SOUND MARK
	`´`: [u8(0x81), 0x4C] // U+00B4 ACUTE ACCENT
	`｀`: [u8(0x81), 0x4D] // U+FF40 FULLWIDTH GRAVE ACCENT
	`¨`: [u8(0x81), 0x4E] // U+00A8 DIAERESIS
	`＾`: [u8(0x81), 0x4F] // U+FF3E FULLWIDTH CIRCUMFLEX ACCENT
	`￣`: [u8(0x81), 0x50] // U+FFE3 FULLWIDTH MACRON
	`＿`: [u8(0x81), 0x51] // U+FF3F FULLWIDTH LOW LINE
	`ヽ`: [u8(0x81), 0x52] // U+30FD KATAKANA ITERATION MARK
	`ヾ`: [u8(0x81), 0x53] // U+30FE KATAKANA VOICED ITERATION MARK
	`ゝ`: [u8(0x81), 0x54] // U+309D HIRAGANA ITERATION MARK
	`ゞ`: [u8(0x81), 0x55] // U+309E HIRAGANA VOICED ITERATION MARK
	`〃`: [u8(0x81), 0x56] // U+3003 DITTO MARK
	`仝`: [u8(0x81), 0x57] // U+4EDD <cjk>
	`々`: [u8(0x81), 0x58] // U+3005 IDEOGRAPHIC ITERATION MARK
	`〆`: [u8(0x81), 0x59] // U+3006 IDEOGRAPHIC CLOSING MARK
	`〇`: [u8(0x81), 0x5A] // U+3007 IDEOGRAPHIC NUMBER ZERO
	`ー`: [u8(0x81), 0x5B] // U+30FC KATAKANA-HIRAGANA PROLONGED SOUND MARK
	`—`: [u8(0x81), 0x5C] // U+2014 EM DASH
	`‐`: [u8(0x81), 0x5D] // U+2010 HYPHEN
	`／`: [u8(0x81), 0x5E] // U+FF0F FULLWIDTH SOLIDUS
	`\\`: [u8(0x81), 0x5F] // U+005C REVERSE SOLIDUS
	`〜`: [u8(0x81), 0x60] // U+301C WAVE DASH
	`‖`: [u8(0x81), 0x61] // U+2016 DOUBLE VERTICAL LINE
	`｜`: [u8(0x81), 0x62] // U+FF5C FULLWIDTH VERTICAL LINE
	`…`: [u8(0x81), 0x63] // U+2026 HORIZONTAL ELLIPSIS
	`‥`: [u8(0x81), 0x64] // U+2025 TWO DOT LEADER
	`‘`: [u8(0x81), 0x65] // U+2018 LEFT SINGLE QUOTATION MARK
	`’`: [u8(0x81), 0x66] // U+2019 RIGHT SINGLE QUOTATION MARK
	`“`: [u8(0x81), 0x67] // U+201C LEFT DOUBLE QUOTATION MARK
	`”`: [u8(0x81), 0x68] // U+201D RIGHT DOUBLE QUOTATION MARK
	`（`: [u8(0x81), 0x69] // U+FF08 FULLWIDTH LEFT PARENTHESIS
	`）`: [u8(0x81), 0x6A] // U+FF09 FULLWIDTH RIGHT PARENTHESIS
	`〔`: [u8(0x81), 0x6B] // U+3014 LEFT TORTOISE SHELL BRACKET
	`〕`: [u8(0x81), 0x6C] // U+3015 RIGHT TORTOISE SHELL BRACKET
	`［`: [u8(0x81), 0x6D] // U+FF3B FULLWIDTH LEFT SQUARE BRACKET
	`］`: [u8(0x81), 0x6E] // U+FF3D FULLWIDTH RIGHT SQUARE BRACKET
	`｛`: [u8(0x81), 0x6F] // U+FF5B FULLWIDTH LEFT CURLY BRACKET
	`｝`: [u8(0x81), 0x70] // U+FF5D FULLWIDTH RIGHT CURLY BRACKET
	`〈`: [u8(0x81), 0x71] // U+3008 LEFT ANGLE BRACKET
	`〉`: [u8(0x81), 0x72] // U+3009 RIGHT ANGLE BRACKET
	`《`: [u8(0x81), 0x73] // U+300A LEFT DOUBLE ANGLE BRACKET
	`》`: [u8(0x81), 0x74] // U+300B RIGHT DOUBLE ANGLE BRACKET
	`「`: [u8(0x81), 0x75] // U+300C LEFT CORNER BRACKET
	`」`: [u8(0x81), 0x76] // U+300D RIGHT CORNER BRACKET
	`『`: [u8(0x81), 0x77] // U+300E LEFT WHITE CORNER BRACKET
	`』`: [u8(0x81), 0x78] // U+300F RIGHT WHITE CORNER BRACKET
	`【`: [u8(0x81), 0x79] // U+3010 LEFT BLACK LENTICULAR BRACKET
	`】`: [u8(0x81), 0x7A] // U+3011 RIGHT BLACK LENTICULAR BRACKET
	`＋`: [u8(0x81), 0x7B] // U+FF0B FULLWIDTH PLUS SIGN
	`−`: [u8(0x81), 0x7C] // U+2212 MINUS SIGN
	`±`: [u8(0x81), 0x7D] // U+00B1 PLUS-MINUS SIGN
	`×`: [u8(0x81), 0x7E] // U+00D7 MULTIPLICATION SIGN
	`÷`: [u8(0x81), 0x80] // U+00F7 DIVISION SIGN
	`＝`: [u8(0x81), 0x81] // U+FF1D FULLWIDTH EQUALS SIGN
	`≠`: [u8(0x81), 0x82] // U+2260 NOT EQUAL TO
	`＜`: [u8(0x81), 0x83] // U+FF1C FULLWIDTH LESS-THAN SIGN
	`＞`: [u8(0x81), 0x84] // U+FF1E FULLWIDTH GREATER-THAN SIGN
	`≦`: [u8(0x81), 0x85] // U+2266 LESS-THAN OVER EQUAL TO
	`≧`: [u8(0x81), 0x86] // U+2267 GREATER-THAN OVER EQUAL TO
	`∞`: [u8(0x81), 0x87] // U+221E INFINITY
	`∴`: [u8(0x81), 0x88] // U+2234 THEREFORE
	`♂`: [u8(0x81), 0x89] // U+2642 MALE SIGN
	`♀`: [u8(0x81), 0x8A] // U+2640 FEMALE SIGN
	`°`: [u8(0x81), 0x8B] // U+00B0 DEGREE SIGN
	`′`: [u8(0x81), 0x8C] // U+2032 PRIME
	`″`: [u8(0x81), 0x8D] // U+2033 DOUBLE PRIME
	`℃`: [u8(0x81), 0x8E] // U+2103 DEGREE CELSIUS
	`￥`: [u8(0x81), 0x8F] // U+FFE5 FULLWIDTH YEN SIGN
	`＄`: [u8(0x81), 0x90] // U+FF04 FULLWIDTH DOLLAR SIGN
	`¢`: [u8(0x81), 0x91] // U+00A2 CENT SIGN
	`£`: [u8(0x81), 0x92] // U+00A3 POUND SIGN
	`％`: [u8(0x81), 0x93] // U+FF05 FULLWIDTH PERCENT SIGN
	`＃`: [u8(0x81), 0x94] // U+FF03 FULLWIDTH NUMBER SIGN
	`＆`: [u8(0x81), 0x95] // U+FF06 FULLWIDTH AMPERSAND
	`＊`: [u8(0x81), 0x96] // U+FF0A FULLWIDTH ASTERISK
	`＠`: [u8(0x81), 0x97] // U+FF20 FULLWIDTH COMMERCIAL AT
	`§`: [u8(0x81), 0x98] // U+00A7 SECTION SIGN
	`☆`: [u8(0x81), 0x99] // U+2606 WHITE STAR
	`★`: [u8(0x81), 0x9A] // U+2605 BLACK STAR
	`○`: [u8(0x81), 0x9B] // U+25CB WHITE CIRCLE
	`●`: [u8(0x81), 0x9C] // U+25CF BLACK CIRCLE
	`◎`: [u8(0x81), 0x9D] // U+25CE BULLSEYE
	`◇`: [u8(0x81), 0x9E] // U+25C7 WHITE DIAMOND
	`◆`: [u8(0x81), 0x9F] // U+25C6 BLACK DIAMOND
	`□`: [u8(0x81), 0xA0] // U+25A1 WHITE SQUARE
	`■`: [u8(0x81), 0xA1] // U+25A0 BLACK SQUARE
	`△`: [u8(0x81), 0xA2] // U+25B3 WHITE UP-POINTING TRIANGLE
	`▲`: [u8(0x81), 0xA3] // U+25B2 BLACK UP-POINTING TRIANGLE
	`▽`: [u8(0x81), 0xA4] // U+25BD WHITE DOWN-POINTING TRIANGLE
	`▼`: [u8(0x81), 0xA5] // U+25BC BLACK DOWN-POINTING TRIANGLE
	`※`: [u8(0x81), 0xA6] // U+203B REFERENCE MARK
	`〒`: [u8(0x81), 0xA7] // U+3012 POSTAL MARK
	`→`: [u8(0x81), 0xA8] // U+2192 RIGHTWARDS ARROW
	`←`: [u8(0x81), 0xA9] // U+2190 LEFTWARDS ARROW
	`↑`: [u8(0x81), 0xAA] // U+2191 UPWARDS ARROW
	`↓`: [u8(0x81), 0xAB] // U+2193 DOWNWARDS ARROW
	`〓`: [u8(0x81), 0xAC] // U+3013 GETA MARK
	`＇`: [u8(0x81), 0xAD] // U+FF07 FULLWIDTH APOSTROPHE
	`＂`: [u8(0x81), 0xAE] // U+FF02 FULLWIDTH QUOTATION MARK
	`－`: [u8(0x81), 0xAF] // U+FF0D FULLWIDTH HYPHEN-MINUS
	`~`: [u8(0x81), 0xB0] // U+007E TILDE
	`〳`: [u8(0x81), 0xB1] // U+3033 VERTICAL KANA REPEAT MARK UPPER HALF
	`〴`: [u8(0x81), 0xB2] // U+3034 VERTICAL KANA REPEAT WITH VOICED SOUND MARK UPPER HALF
	`〵`: [u8(0x81), 0xB3] // U+3035 VERTICAL KANA REPEAT MARK LOWER HALF
	`〻`: [u8(0x81), 0xB4] // U+303B VERTICAL IDEOGRAPHIC ITERATION MARK
	`〼`: [u8(0x81), 0xB5] // U+303C MASU MARK
	`ヿ`: [u8(0x81), 0xB6] // U+30FF KATAKANA DIGRAPH KOTO
	`ゟ`: [u8(0x81), 0xB7] // U+309F HIRAGANA DIGRAPH YORI
	`∈`: [u8(0x81), 0xB8] // U+2208 ELEMENT OF
	`∋`: [u8(0x81), 0xB9] // U+220B CONTAINS AS MEMBER
	`⊆`: [u8(0x81), 0xBA] // U+2286 SUBSET OF OR EQUAL TO
	`⊇`: [u8(0x81), 0xBB] // U+2287 SUPERSET OF OR EQUAL TO
	`⊂`: [u8(0x81), 0xBC] // U+2282 SUBSET OF
	`⊃`: [u8(0x81), 0xBD] // U+2283 SUPERSET OF
	`∪`: [u8(0x81), 0xBE] // U+222A UNION
	`∩`: [u8(0x81), 0xBF] // U+2229 INTERSECTION
	`⊄`: [u8(0x81), 0xC0] // U+2284 NOT A SUBSET OF
	`⊅`: [u8(0x81), 0xC1] // U+2285 NOT A SUPERSET OF
	`⊊`: [u8(0x81), 0xC2] // U+228A SUBSET OF WITH NOT EQUAL TO
	`⊋`: [u8(0x81), 0xC3] // U+228B SUPERSET OF WITH NOT EQUAL TO
	`∉`: [u8(0x81), 0xC4] // U+2209 NOT AN ELEMENT OF
	`∅`: [u8(0x81), 0xC5] // U+2205 EMPTY SET
	`⌅`: [u8(0x81), 0xC6] // U+2305 PROJECTIVE
	`⌆`: [u8(0x81), 0xC7] // U+2306 PERSPECTIVE
	`∧`: [u8(0x81), 0xC8] // U+2227 LOGICAL AND
	`∨`: [u8(0x81), 0xC9] // U+2228 LOGICAL OR
	`¬`: [u8(0x81), 0xCA] // U+00AC NOT SIGN
	`⇒`: [u8(0x81), 0xCB] // U+21D2 RIGHTWARDS DOUBLE ARROW
	`⇔`: [u8(0x81), 0xCC] // U+21D4 LEFT RIGHT DOUBLE ARROW
	`∀`: [u8(0x81), 0xCD] // U+2200 FOR ALL
	`∃`: [u8(0x81), 0xCE] // U+2203 THERE EXISTS
	`⊕`: [u8(0x81), 0xCF] // U+2295 CIRCLED PLUS
	`⊖`: [u8(0x81), 0xD0] // U+2296 CIRCLED MINUS
	`⊗`: [u8(0x81), 0xD1] // U+2297 CIRCLED TIMES
	`∥`: [u8(0x81), 0xD2] // U+2225 PARALLEL TO
	`∦`: [u8(0x81), 0xD3] // U+2226 NOT PARALLEL TO
	`｟`: [u8(0x81), 0xD4] // U+FF5F FULLWIDTH LEFT WHITE PARENTHESIS
	`｠`: [u8(0x81), 0xD5] // U+FF60 FULLWIDTH RIGHT WHITE PARENTHESIS
	`〘`: [u8(0x81), 0xD6] // U+3018 LEFT WHITE TORTOISE SHELL BRACKET
	`〙`: [u8(0x81), 0xD7] // U+3019 RIGHT WHITE TORTOISE SHELL BRACKET
	`〖`: [u8(0x81), 0xD8] // U+3016 LEFT WHITE LENTICULAR BRACKET
	`〗`: [u8(0x81), 0xD9] // U+3017 RIGHT WHITE LENTICULAR BRACKET
	`∠`: [u8(0x81), 0xDA] // U+2220 ANGLE
	`⊥`: [u8(0x81), 0xDB] // U+22A5 UP TACK
	`⌒`: [u8(0x81), 0xDC] // U+2312 ARC
	`∂`: [u8(0x81), 0xDD] // U+2202 PARTIAL DIFFERENTIAL
	`∇`: [u8(0x81), 0xDE] // U+2207 NABLA
	`≡`: [u8(0x81), 0xDF] // U+2261 IDENTICAL TO
	`≒`: [u8(0x81), 0xE0] // U+2252 APPROXIMATELY EQUAL TO OR THE IMAGE OF
	`≪`: [u8(0x81), 0xE1] // U+226A MUCH LESS-THAN
	`≫`: [u8(0x81), 0xE2] // U+226B MUCH GREATER-THAN
	`√`: [u8(0x81), 0xE3] // U+221A SQUARE ROOT
	`∽`: [u8(0x81), 0xE4] // U+223D REVERSED TILDE
	`∝`: [u8(0x81), 0xE5] // U+221D PROPORTIONAL TO
	`∵`: [u8(0x81), 0xE6] // U+2235 BECAUSE
	`∫`: [u8(0x81), 0xE7] // U+222B INTEGRAL
	`∬`: [u8(0x81), 0xE8] // U+222C DOUBLE INTEGRAL
	`≢`: [u8(0x81), 0xE9] // U+2262 NOT IDENTICAL TO
	`≃`: [u8(0x81), 0xEA] // U+2243 ASYMPTOTICALLY EQUAL TO
	`≅`: [u8(0x81), 0xEB] // U+2245 APPROXIMATELY EQUAL TO
	`≈`: [u8(0x81), 0xEC] // U+2248 ALMOST EQUAL TO
	`≶`: [u8(0x81), 0xED] // U+2276 LESS-THAN OR GREATER-THAN
	`≷`: [u8(0x81), 0xEE] // U+2277 GREATER-THAN OR LESS-THAN
	`↔`: [u8(0x81), 0xEF] // U+2194 LEFT RIGHT ARROW
	`Å`: [u8(0x81), 0xF0] // U+212B ANGSTROM SIGN
	`‰`: [u8(0x81), 0xF1] // U+2030 PER MILLE SIGN
	`♯`: [u8(0x81), 0xF2] // U+266F MUSIC SHARP SIGN
	`♭`: [u8(0x81), 0xF3] // U+266D MUSIC FLAT SIGN
	`♪`: [u8(0x81), 0xF4] // U+266A EIGHTH NOTE
	`†`: [u8(0x81), 0xF5] // U+2020 DAGGER
	`‡`: [u8(0x81), 0xF6] // U+2021 DOUBLE DAGGER
	`¶`: [u8(0x81), 0xF7] // U+00B6 PILCROW SIGN
	`♮`: [u8(0x81), 0xF8] // U+266E MUSIC NATURAL SIGN
	`♫`: [u8(0x81), 0xF9] // U+266B BEAMED EIGHTH NOTES
	`♬`: [u8(0x81), 0xFA] // U+266C BEAMED SIXTEENTH NOTES
	`♩`: [u8(0x81), 0xFB] // U+2669 QUARTER NOTE
	`◯`: [u8(0x81), 0xFC] // U+25EF LARGE CIRCLE
	`▷`: [u8(0x82), 0x40] // U+25B7 WHITE RIGHT-POINTING TRIANGLE
	`▶`: [u8(0x82), 0x41] // U+25B6 BLACK RIGHT-POINTING TRIANGLE
	`◁`: [u8(0x82), 0x42] // U+25C1 WHITE LEFT-POINTING TRIANGLE
	`◀`: [u8(0x82), 0x43] // U+25C0 BLACK LEFT-POINTING TRIANGLE
	`↗`: [u8(0x82), 0x44] // U+2197 NORTH EAST ARROW
	`↘`: [u8(0x82), 0x45] // U+2198 SOUTH EAST ARROW
	`↖`: [u8(0x82), 0x46] // U+2196 NORTH WEST ARROW
	`↙`: [u8(0x82), 0x47] // U+2199 SOUTH WEST ARROW
	`⇄`: [u8(0x82), 0x48] // U+21C4 RIGHTWARDS ARROW OVER LEFTWARDS ARROW
	`⇨`: [u8(0x82), 0x49] // U+21E8 RIGHTWARDS WHITE ARROW
	`⇦`: [u8(0x82), 0x4A] // U+21E6 LEFTWARDS WHITE ARROW
	`⇧`: [u8(0x82), 0x4B] // U+21E7 UPWARDS WHITE ARROW
	`⇩`: [u8(0x82), 0x4C] // U+21E9 DOWNWARDS WHITE ARROW
	`⤴`: [u8(0x82), 0x4D] // U+2934 ARROW POINTING RIGHTWARDS THEN CURVING UPWARDS
	`⤵`: [u8(0x82), 0x4E] // U+2935 ARROW POINTING RIGHTWARDS THEN CURVING DOWNWARDS
	`０`: [u8(0x82), 0x4F] // U+FF10 FULLWIDTH DIGIT ZERO
	`１`: [u8(0x82), 0x50] // U+FF11 FULLWIDTH DIGIT ONE
	`２`: [u8(0x82), 0x51] // U+FF12 FULLWIDTH DIGIT TWO
	`３`: [u8(0x82), 0x52] // U+FF13 FULLWIDTH DIGIT THREE
	`４`: [u8(0x82), 0x53] // U+FF14 FULLWIDTH DIGIT FOUR
	`５`: [u8(0x82), 0x54] // U+FF15 FULLWIDTH DIGIT FIVE
	`６`: [u8(0x82), 0x55] // U+FF16 FULLWIDTH DIGIT SIX
	`７`: [u8(0x82), 0x56] // U+FF17 FULLWIDTH DIGIT SEVEN
	`８`: [u8(0x82), 0x57] // U+FF18 FULLWIDTH DIGIT EIGHT
	`９`: [u8(0x82), 0x58] // U+FF19 FULLWIDTH DIGIT NINE
	`⦿`: [u8(0x82), 0x59] // U+29BF CIRCLED BULLET
	`◉`: [u8(0x82), 0x5A] // U+25C9 FISHEYE
	`〽`: [u8(0x82), 0x5B] // U+303D PART ALTERNATION MARK
	`﹆`: [u8(0x82), 0x5C] // U+FE46 WHITE SESAME DOT
	`﹅`: [u8(0x82), 0x5D] // U+FE45 SESAME DOT
	`◦`: [u8(0x82), 0x5E] // U+25E6 WHITE BULLET
	`•`: [u8(0x82), 0x5F] // U+2022 BULLET
	`Ａ`: [u8(0x82), 0x60] // U+FF21 FULLWIDTH LATIN CAPITAL LETTER A
	`Ｂ`: [u8(0x82), 0x61] // U+FF22 FULLWIDTH LATIN CAPITAL LETTER B
	`Ｃ`: [u8(0x82), 0x62] // U+FF23 FULLWIDTH LATIN CAPITAL LETTER C
	`Ｄ`: [u8(0x82), 0x63] // U+FF24 FULLWIDTH LATIN CAPITAL LETTER D
	`Ｅ`: [u8(0x82), 0x64] // U+FF25 FULLWIDTH LATIN CAPITAL LETTER E
	`Ｆ`: [u8(0x82), 0x65] // U+FF26 FULLWIDTH LATIN CAPITAL LETTER F
	`Ｇ`: [u8(0x82), 0x66] // U+FF27 FULLWIDTH LATIN CAPITAL LETTER G
	`Ｈ`: [u8(0x82), 0x67] // U+FF28 FULLWIDTH LATIN CAPITAL LETTER H
	`Ｉ`: [u8(0x82), 0x68] // U+FF29 FULLWIDTH LATIN CAPITAL LETTER I
	`Ｊ`: [u8(0x82), 0x69] // U+FF2A FULLWIDTH LATIN CAPITAL LETTER J
	`Ｋ`: [u8(0x82), 0x6A] // U+FF2B FULLWIDTH LATIN CAPITAL LETTER K
	`Ｌ`: [u8(0x82), 0x6B] // U+FF2C FULLWIDTH LATIN CAPITAL LETTER L
	`Ｍ`: [u8(0x82), 0x6C] // U+FF2D FULLWIDTH LATIN CAPITAL LETTER M
	`Ｎ`: [u8(0x82), 0x6D] // U+FF2E FULLWIDTH LATIN CAPITAL LETTER N
	`Ｏ`: [u8(0x82), 0x6E] // U+FF2F FULLWIDTH LATIN CAPITAL LETTER O
	`Ｐ`: [u8(0x82), 0x6F] // U+FF30 FULLWIDTH LATIN CAPITAL LETTER P
	`Ｑ`: [u8(0x82), 0x70] // U+FF31 FULLWIDTH LATIN CAPITAL LETTER Q
	`Ｒ`: [u8(0x82), 0x71] // U+FF32 FULLWIDTH LATIN CAPITAL LETTER R
	`Ｓ`: [u8(0x82), 0x72] // U+FF33 FULLWIDTH LATIN CAPITAL LETTER S
	`Ｔ`: [u8(0x82), 0x73] // U+FF34 FULLWIDTH LATIN CAPITAL LETTER T
	`Ｕ`: [u8(0x82), 0x74] // U+FF35 FULLWIDTH LATIN CAPITAL LETTER U
	`Ｖ`: [u8(0x82), 0x75] // U+FF36 FULLWIDTH LATIN CAPITAL LETTER V
	`Ｗ`: [u8(0x82), 0x76] // U+FF37 FULLWIDTH LATIN CAPITAL LETTER W
	`Ｘ`: [u8(0x82), 0x77] // U+FF38 FULLWIDTH LATIN CAPITAL LETTER X
	`Ｙ`: [u8(0x82), 0x78] // U+FF39 FULLWIDTH LATIN CAPITAL LETTER Y
	`Ｚ`: [u8(0x82), 0x79] // U+FF3A FULLWIDTH LATIN CAPITAL LETTER Z
	`∓`: [u8(0x82), 0x7A] // U+2213 MINUS-OR-PLUS SIGN
	`ℵ`: [u8(0x82), 0x7B] // U+2135 ALEF SYMBOL
	`ℏ`: [u8(0x82), 0x7C] // U+210F PLANCK CONSTANT OVER TWO PI
	`㏋`: [u8(0x82), 0x7D] // U+33CB SQUARE HP
	`ℓ`: [u8(0x82), 0x7E] // U+2113 SCRIPT SMALL L
	`℧`: [u8(0x82), 0x80] // U+2127 INVERTED OHM SIGN
	`ａ`: [u8(0x82), 0x81] // U+FF41 FULLWIDTH LATIN SMALL LETTER A
	`ｂ`: [u8(0x82), 0x82] // U+FF42 FULLWIDTH LATIN SMALL LETTER B
	`ｃ`: [u8(0x82), 0x83] // U+FF43 FULLWIDTH LATIN SMALL LETTER C
	`ｄ`: [u8(0x82), 0x84] // U+FF44 FULLWIDTH LATIN SMALL LETTER D
	`ｅ`: [u8(0x82), 0x85] // U+FF45 FULLWIDTH LATIN SMALL LETTER E
	`ｆ`: [u8(0x82), 0x86] // U+FF46 FULLWIDTH LATIN SMALL LETTER F
	`ｇ`: [u8(0x82), 0x87] // U+FF47 FULLWIDTH LATIN SMALL LETTER G
	`ｈ`: [u8(0x82), 0x88] // U+FF48 FULLWIDTH LATIN SMALL LETTER H
	`ｉ`: [u8(0x82), 0x89] // U+FF49 FULLWIDTH LATIN SMALL LETTER I
	`ｊ`: [u8(0x82), 0x8A] // U+FF4A FULLWIDTH LATIN SMALL LETTER J
	`ｋ`: [u8(0x82), 0x8B] // U+FF4B FULLWIDTH LATIN SMALL LETTER K
	`ｌ`: [u8(0x82), 0x8C] // U+FF4C FULLWIDTH LATIN SMALL LETTER L
	`ｍ`: [u8(0x82), 0x8D] // U+FF4D FULLWIDTH LATIN SMALL LETTER M
	`ｎ`: [u8(0x82), 0x8E] // U+FF4E FULLWIDTH LATIN SMALL LETTER N
	`ｏ`: [u8(0x82), 0x8F] // U+FF4F FULLWIDTH LATIN SMALL LETTER O
	`ｐ`: [u8(0x82), 0x90] // U+FF50 FULLWIDTH LATIN SMALL LETTER P
	`ｑ`: [u8(0x82), 0x91] // U+FF51 FULLWIDTH LATIN SMALL LETTER Q
	`ｒ`: [u8(0x82), 0x92] // U+FF52 FULLWIDTH LATIN SMALL LETTER R
	`ｓ`: [u8(0x82), 0x93] // U+FF53 FULLWIDTH LATIN SMALL LETTER S
	`ｔ`: [u8(0x82), 0x94] // U+FF54 FULLWIDTH LATIN SMALL LETTER T
	`ｕ`: [u8(0x82), 0x95] // U+FF55 FULLWIDTH LATIN SMALL LETTER U
	`ｖ`: [u8(0x82), 0x96] // U+FF56 FULLWIDTH LATIN SMALL LETTER V
	`ｗ`: [u8(0x82), 0x97] // U+FF57 FULLWIDTH LATIN SMALL LETTER W
	`ｘ`: [u8(0x82), 0x98] // U+FF58 FULLWIDTH LATIN SMALL LETTER X
	`ｙ`: [u8(0x82), 0x99] // U+FF59 FULLWIDTH LATIN SMALL LETTER Y
	`ｚ`: [u8(0x82), 0x9A] // U+FF5A FULLWIDTH LATIN SMALL LETTER Z
	`゠`: [u8(0x82), 0x9B] // U+30A0 KATAKANA-HIRAGANA DOUBLE HYPHEN
	`–`: [u8(0x82), 0x9C] // U+2013 EN DASH
	`⧺`: [u8(0x82), 0x9D] // U+29FA DOUBLE PLUS
	`⧻`: [u8(0x82), 0x9E] // U+29FB TRIPLE PLUS
	`ぁ`: [u8(0x82), 0x9F] // U+3041 HIRAGANA LETTER SMALL A
	`あ`: [u8(0x82), 0xA0] // U+3042 HIRAGANA LETTER A
	`ぃ`: [u8(0x82), 0xA1] // U+3043 HIRAGANA LETTER SMALL I
	`い`: [u8(0x82), 0xA2] // U+3044 HIRAGANA LETTER I
	`ぅ`: [u8(0x82), 0xA3] // U+3045 HIRAGANA LETTER SMALL U
	`う`: [u8(0x82), 0xA4] // U+3046 HIRAGANA LETTER U
	`ぇ`: [u8(0x82), 0xA5] // U+3047 HIRAGANA LETTER SMALL E
	`え`: [u8(0x82), 0xA6] // U+3048 HIRAGANA LETTER E
	`ぉ`: [u8(0x82), 0xA7] // U+3049 HIRAGANA LETTER SMALL O
	`お`: [u8(0x82), 0xA8] // U+304A HIRAGANA LETTER O
	`か`: [u8(0x82), 0xA9] // U+304B HIRAGANA LETTER KA
	`が`: [u8(0x82), 0xAA] // U+304C HIRAGANA LETTER GA
	`き`: [u8(0x82), 0xAB] // U+304D HIRAGANA LETTER KI
	`ぎ`: [u8(0x82), 0xAC] // U+304E HIRAGANA LETTER GI
	`く`: [u8(0x82), 0xAD] // U+304F HIRAGANA LETTER KU
	`ぐ`: [u8(0x82), 0xAE] // U+3050 HIRAGANA LETTER GU
	`け`: [u8(0x82), 0xAF] // U+3051 HIRAGANA LETTER KE
	`げ`: [u8(0x82), 0xB0] // U+3052 HIRAGANA LETTER GE
	`こ`: [u8(0x82), 0xB1] // U+3053 HIRAGANA LETTER KO
	`ご`: [u8(0x82), 0xB2] // U+3054 HIRAGANA LETTER GO
	`さ`: [u8(0x82), 0xB3] // U+3055 HIRAGANA LETTER SA
	`ざ`: [u8(0x82), 0xB4] // U+3056 HIRAGANA LETTER ZA
	`し`: [u8(0x82), 0xB5] // U+3057 HIRAGANA LETTER SI
	`じ`: [u8(0x82), 0xB6] // U+3058 HIRAGANA LETTER ZI
	`す`: [u8(0x82), 0xB7] // U+3059 HIRAGANA LETTER SU
	`ず`: [u8(0x82), 0xB8] // U+305A HIRAGANA LETTER ZU
	`せ`: [u8(0x82), 0xB9] // U+305B HIRAGANA LETTER SE
	`ぜ`: [u8(0x82), 0xBA] // U+305C HIRAGANA LETTER ZE
	`そ`: [u8(0x82), 0xBB] // U+305D HIRAGANA LETTER SO
	`ぞ`: [u8(0x82), 0xBC] // U+305E HIRAGANA LETTER ZO
	`た`: [u8(0x82), 0xBD] // U+305F HIRAGANA LETTER TA
	`だ`: [u8(0x82), 0xBE] // U+3060 HIRAGANA LETTER DA
	`ち`: [u8(0x82), 0xBF] // U+3061 HIRAGANA LETTER TI
	`ぢ`: [u8(0x82), 0xC0] // U+3062 HIRAGANA LETTER DI
	`っ`: [u8(0x82), 0xC1] // U+3063 HIRAGANA LETTER SMALL TU
	`つ`: [u8(0x82), 0xC2] // U+3064 HIRAGANA LETTER TU
	`づ`: [u8(0x82), 0xC3] // U+3065 HIRAGANA LETTER DU
	`て`: [u8(0x82), 0xC4] // U+3066 HIRAGANA LETTER TE
	`で`: [u8(0x82), 0xC5] // U+3067 HIRAGANA LETTER DE
	`と`: [u8(0x82), 0xC6] // U+3068 HIRAGANA LETTER TO
	`ど`: [u8(0x82), 0xC7] // U+3069 HIRAGANA LETTER DO
	`な`: [u8(0x82), 0xC8] // U+306A HIRAGANA LETTER NA
	`に`: [u8(0x82), 0xC9] // U+306B HIRAGANA LETTER NI
	`ぬ`: [u8(0x82), 0xCA] // U+306C HIRAGANA LETTER NU
	`ね`: [u8(0x82), 0xCB] // U+306D HIRAGANA LETTER NE
	`の`: [u8(0x82), 0xCC] // U+306E HIRAGANA LETTER NO
	`は`: [u8(0x82), 0xCD] // U+306F HIRAGANA LETTER HA
	`ば`: [u8(0x82), 0xCE] // U+3070 HIRAGANA LETTER BA
	`ぱ`: [u8(0x82), 0xCF] // U+3071 HIRAGANA LETTER PA
	`ひ`: [u8(0x82), 0xD0] // U+3072 HIRAGANA LETTER HI
	`び`: [u8(0x82), 0xD1] // U+3073 HIRAGANA LETTER BI
	`ぴ`: [u8(0x82), 0xD2] // U+3074 HIRAGANA LETTER PI
	`ふ`: [u8(0x82), 0xD3] // U+3075 HIRAGANA LETTER HU
	`ぶ`: [u8(0x82), 0xD4] // U+3076 HIRAGANA LETTER BU
	`ぷ`: [u8(0x82), 0xD5] // U+3077 HIRAGANA LETTER PU
	`へ`: [u8(0x82), 0xD6] // U+3078 HIRAGANA LETTER HE
	`べ`: [u8(0x82), 0xD7] // U+3079 HIRAGANA LETTER BE
	`ぺ`: [u8(0x82), 0xD8] // U+307A HIRAGANA LETTER PE
	`ほ`: [u8(0x82), 0xD9] // U+307B HIRAGANA LETTER HO
	`ぼ`: [u8(0x82), 0xDA] // U+307C HIRAGANA LETTER BO
	`ぽ`: [u8(0x82), 0xDB] // U+307D HIRAGANA LETTER PO
	`ま`: [u8(0x82), 0xDC] // U+307E HIRAGANA LETTER MA
	`み`: [u8(0x82), 0xDD] // U+307F HIRAGANA LETTER MI
	`む`: [u8(0x82), 0xDE] // U+3080 HIRAGANA LETTER MU
	`め`: [u8(0x82), 0xDF] // U+3081 HIRAGANA LETTER ME
	`も`: [u8(0x82), 0xE0] // U+3082 HIRAGANA LETTER MO
	`ゃ`: [u8(0x82), 0xE1] // U+3083 HIRAGANA LETTER SMALL YA
	`や`: [u8(0x82), 0xE2] // U+3084 HIRAGANA LETTER YA
	`ゅ`: [u8(0x82), 0xE3] // U+3085 HIRAGANA LETTER SMALL YU
	`ゆ`: [u8(0x82), 0xE4] // U+3086 HIRAGANA LETTER YU
	`ょ`: [u8(0x82), 0xE5] // U+3087 HIRAGANA LETTER SMALL YO
	`よ`: [u8(0x82), 0xE6] // U+3088 HIRAGANA LETTER YO
	`ら`: [u8(0x82), 0xE7] // U+3089 HIRAGANA LETTER RA
	`り`: [u8(0x82), 0xE8] // U+308A HIRAGANA LETTER RI
	`る`: [u8(0x82), 0xE9] // U+308B HIRAGANA LETTER RU
	`れ`: [u8(0x82), 0xEA] // U+308C HIRAGANA LETTER RE
	`ろ`: [u8(0x82), 0xEB] // U+308D HIRAGANA LETTER RO
	`ゎ`: [u8(0x82), 0xEC] // U+308E HIRAGANA LETTER SMALL WA
	`わ`: [u8(0x82), 0xED] // U+308F HIRAGANA LETTER WA
	`ゐ`: [u8(0x82), 0xEE] // U+3090 HIRAGANA LETTER WI
	`ゑ`: [u8(0x82), 0xEF] // U+3091 HIRAGANA LETTER WE
	`を`: [u8(0x82), 0xF0] // U+3092 HIRAGANA LETTER WO
	`ん`: [u8(0x82), 0xF1] // U+3093 HIRAGANA LETTER N
	`ゔ`: [u8(0x82), 0xF2] // U+3094 HIRAGANA LETTER VU
	`ゕ`: [u8(0x82), 0xF3] // U+3095 HIRAGANA LETTER SMALL KA
	`ゖ`: [u8(0x82), 0xF4] // U+3096 HIRAGANA LETTER SMALL KE
	`ァ`: [u8(0x83), 0x40] // U+30A1 KATAKANA LETTER SMALL A
	`ア`: [u8(0x83), 0x41] // U+30A2 KATAKANA LETTER A
	`ィ`: [u8(0x83), 0x42] // U+30A3 KATAKANA LETTER SMALL I
	`イ`: [u8(0x83), 0x43] // U+30A4 KATAKANA LETTER I
	`ゥ`: [u8(0x83), 0x44] // U+30A5 KATAKANA LETTER SMALL U
	`ウ`: [u8(0x83), 0x45] // U+30A6 KATAKANA LETTER U
	`ェ`: [u8(0x83), 0x46] // U+30A7 KATAKANA LETTER SMALL E
	`エ`: [u8(0x83), 0x47] // U+30A8 KATAKANA LETTER E
	`ォ`: [u8(0x83), 0x48] // U+30A9 KATAKANA LETTER SMALL O
	`オ`: [u8(0x83), 0x49] // U+30AA KATAKANA LETTER O
	`カ`: [u8(0x83), 0x4A] // U+30AB KATAKANA LETTER KA
	`ガ`: [u8(0x83), 0x4B] // U+30AC KATAKANA LETTER GA
	`キ`: [u8(0x83), 0x4C] // U+30AD KATAKANA LETTER KI
	`ギ`: [u8(0x83), 0x4D] // U+30AE KATAKANA LETTER GI
	`ク`: [u8(0x83), 0x4E] // U+30AF KATAKANA LETTER KU
	`グ`: [u8(0x83), 0x4F] // U+30B0 KATAKANA LETTER GU
	`ケ`: [u8(0x83), 0x50] // U+30B1 KATAKANA LETTER KE
	`ゲ`: [u8(0x83), 0x51] // U+30B2 KATAKANA LETTER GE
	`コ`: [u8(0x83), 0x52] // U+30B3 KATAKANA LETTER KO
	`ゴ`: [u8(0x83), 0x53] // U+30B4 KATAKANA LETTER GO
	`サ`: [u8(0x83), 0x54] // U+30B5 KATAKANA LETTER SA
	`ザ`: [u8(0x83), 0x55] // U+30B6 KATAKANA LETTER ZA
	`シ`: [u8(0x83), 0x56] // U+30B7 KATAKANA LETTER SI
	`ジ`: [u8(0x83), 0x57] // U+30B8 KATAKANA LETTER ZI
	`ス`: [u8(0x83), 0x58] // U+30B9 KATAKANA LETTER SU
	`ズ`: [u8(0x83), 0x59] // U+30BA KATAKANA LETTER ZU
	`セ`: [u8(0x83), 0x5A] // U+30BB KATAKANA LETTER SE
	`ゼ`: [u8(0x83), 0x5B] // U+30BC KATAKANA LETTER ZE
	`ソ`: [u8(0x83), 0x5C] // U+30BD KATAKANA LETTER SO
	`ゾ`: [u8(0x83), 0x5D] // U+30BE KATAKANA LETTER ZO
	`タ`: [u8(0x83), 0x5E] // U+30BF KATAKANA LETTER TA
	`ダ`: [u8(0x83), 0x5F] // U+30C0 KATAKANA LETTER DA
	`チ`: [u8(0x83), 0x60] // U+30C1 KATAKANA LETTER TI
	`ヂ`: [u8(0x83), 0x61] // U+30C2 KATAKANA LETTER DI
	`ッ`: [u8(0x83), 0x62] // U+30C3 KATAKANA LETTER SMALL TU
	`ツ`: [u8(0x83), 0x63] // U+30C4 KATAKANA LETTER TU
	`ヅ`: [u8(0x83), 0x64] // U+30C5 KATAKANA LETTER DU
	`テ`: [u8(0x83), 0x65] // U+30C6 KATAKANA LETTER TE
	`デ`: [u8(0x83), 0x66] // U+30C7 KATAKANA LETTER DE
	`ト`: [u8(0x83), 0x67] // U+30C8 KATAKANA LETTER TO
	`ド`: [u8(0x83), 0x68] // U+30C9 KATAKANA LETTER DO
	`ナ`: [u8(0x83), 0x69] // U+30CA KATAKANA LETTER NA
	`ニ`: [u8(0x83), 0x6A] // U+30CB KATAKANA LETTER NI
	`ヌ`: [u8(0x83), 0x6B] // U+30CC KATAKANA LETTER NU
	`ネ`: [u8(0x83), 0x6C] // U+30CD KATAKANA LETTER NE
	`ノ`: [u8(0x83), 0x6D] // U+30CE KATAKANA LETTER NO
	`ハ`: [u8(0x83), 0x6E] // U+30CF KATAKANA LETTER HA
	`バ`: [u8(0x83), 0x6F] // U+30D0 KATAKANA LETTER BA
	`パ`: [u8(0x83), 0x70] // U+30D1 KATAKANA LETTER PA
	`ヒ`: [u8(0x83), 0x71] // U+30D2 KATAKANA LETTER HI
	`ビ`: [u8(0x83), 0x72] // U+30D3 KATAKANA LETTER BI
	`ピ`: [u8(0x83), 0x73] // U+30D4 KATAKANA LETTER PI
	`フ`: [u8(0x83), 0x74] // U+30D5 KATAKANA LETTER HU
	`ブ`: [u8(0x83), 0x75] // U+30D6 KATAKANA LETTER BU
	`プ`: [u8(0x83), 0x76] // U+30D7 KATAKANA LETTER PU
	`ヘ`: [u8(0x83), 0x77] // U+30D8 KATAKANA LETTER HE
	`ベ`: [u8(0x83), 0x78] // U+30D9 KATAKANA LETTER BE
	`ペ`: [u8(0x83), 0x79] // U+30DA KATAKANA LETTER PE
	`ホ`: [u8(0x83), 0x7A] // U+30DB KATAKANA LETTER HO
	`ボ`: [u8(0x83), 0x7B] // U+30DC KATAKANA LETTER BO
	`ポ`: [u8(0x83), 0x7C] // U+30DD KATAKANA LETTER PO
	`マ`: [u8(0x83), 0x7D] // U+30DE KATAKANA LETTER MA
	`ミ`: [u8(0x83), 0x7E] // U+30DF KATAKANA LETTER MI
	`ム`: [u8(0x83), 0x80] // U+30E0 KATAKANA LETTER MU
	`メ`: [u8(0x83), 0x81] // U+30E1 KATAKANA LETTER ME
	`モ`: [u8(0x83), 0x82] // U+30E2 KATAKANA LETTER MO
	`ャ`: [u8(0x83), 0x83] // U+30E3 KATAKANA LETTER SMALL YA
	`ヤ`: [u8(0x83), 0x84] // U+30E4 KATAKANA LETTER YA
	`ュ`: [u8(0x83), 0x85] // U+30E5 KATAKANA LETTER SMALL YU
	`ユ`: [u8(0x83), 0x86] // U+30E6 KATAKANA LETTER YU
	`ョ`: [u8(0x83), 0x87] // U+30E7 KATAKANA LETTER SMALL YO
	`ヨ`: [u8(0x83), 0x88] // U+30E8 KATAKANA LETTER YO
	`ラ`: [u8(0x83), 0x89] // U+30E9 KATAKANA LETTER RA
	`リ`: [u8(0x83), 0x8A] // U+30EA KATAKANA LETTER RI
	`ル`: [u8(0x83), 0x8B] // U+30EB KATAKANA LETTER RU
	`レ`: [u8(0x83), 0x8C] // U+30EC KATAKANA LETTER RE
	`ロ`: [u8(0x83), 0x8D] // U+30ED KATAKANA LETTER RO
	`ヮ`: [u8(0x83), 0x8E] // U+30EE KATAKANA LETTER SMALL WA
	`ワ`: [u8(0x83), 0x8F] // U+30EF KATAKANA LETTER WA
	`ヰ`: [u8(0x83), 0x90] // U+30F0 KATAKANA LETTER WI
	`ヱ`: [u8(0x83), 0x91] // U+30F1 KATAKANA LETTER WE
	`ヲ`: [u8(0x83), 0x92] // U+30F2 KATAKANA LETTER WO
	`ン`: [u8(0x83), 0x93] // U+30F3 KATAKANA LETTER N
	`ヴ`: [u8(0x83), 0x94] // U+30F4 KATAKANA LETTER VU
	`ヵ`: [u8(0x83), 0x95] // U+30F5 KATAKANA LETTER SMALL KA
	`ヶ`: [u8(0x83), 0x96] // U+30F6 KATAKANA LETTER SMALL KE
	`Α`: [u8(0x83), 0x9F] // U+0391 GREEK CAPITAL LETTER ALPHA
	`Β`: [u8(0x83), 0xA0] // U+0392 GREEK CAPITAL LETTER BETA
	`Γ`: [u8(0x83), 0xA1] // U+0393 GREEK CAPITAL LETTER GAMMA
	`Δ`: [u8(0x83), 0xA2] // U+0394 GREEK CAPITAL LETTER DELTA
	`Ε`: [u8(0x83), 0xA3] // U+0395 GREEK CAPITAL LETTER EPSILON
	`Ζ`: [u8(0x83), 0xA4] // U+0396 GREEK CAPITAL LETTER ZETA
	`Η`: [u8(0x83), 0xA5] // U+0397 GREEK CAPITAL LETTER ETA
	`Θ`: [u8(0x83), 0xA6] // U+0398 GREEK CAPITAL LETTER THETA
	`Ι`: [u8(0x83), 0xA7] // U+0399 GREEK CAPITAL LETTER IOTA
	`Κ`: [u8(0x83), 0xA8] // U+039A GREEK CAPITAL LETTER KAPPA
	`Λ`: [u8(0x83), 0xA9] // U+039B GREEK CAPITAL LETTER LAMDA
	`Μ`: [u8(0x83), 0xAA] // U+039C GREEK CAPITAL LETTER MU
	`Ν`: [u8(0x83), 0xAB] // U+039D GREEK CAPITAL LETTER NU
	`Ξ`: [u8(0x83), 0xAC] // U+039E GREEK CAPITAL LETTER XI
	`Ο`: [u8(0x83), 0xAD] // U+039F GREEK CAPITAL LETTER OMICRON
	`Π`: [u8(0x83), 0xAE] // U+03A0 GREEK CAPITAL LETTER PI
	`Ρ`: [u8(0x83), 0xAF] // U+03A1 GREEK CAPITAL LETTER RHO
	`Σ`: [u8(0x83), 0xB0] // U+03A3 GREEK CAPITAL LETTER SIGMA
	`Τ`: [u8(0x83), 0xB1] // U+03A4 GREEK CAPITAL LETTER TAU
	`Υ`: [u8(0x83), 0xB2] // U+03A5 GREEK CAPITAL LETTER UPSILON
	`Φ`: [u8(0x83), 0xB3] // U+03A6 GREEK CAPITAL LETTER PHI
	`Χ`: [u8(0x83), 0xB4] // U+03A7 GREEK CAPITAL LETTER CHI
	`Ψ`: [u8(0x83), 0xB5] // U+03A8 GREEK CAPITAL LETTER PSI
	`Ω`: [u8(0x83), 0xB6] // U+03A9 GREEK CAPITAL LETTER OMEGA
	`♤`: [u8(0x83), 0xB7] // U+2664 WHITE SPADE SUIT
	`♠`: [u8(0x83), 0xB8] // U+2660 BLACK SPADE SUIT
	`♢`: [u8(0x83), 0xB9] // U+2662 WHITE DIAMOND SUIT
	`♦`: [u8(0x83), 0xBA] // U+2666 BLACK DIAMOND SUIT
	`♡`: [u8(0x83), 0xBB] // U+2661 WHITE HEART SUIT
	`♥`: [u8(0x83), 0xBC] // U+2665 BLACK HEART SUIT
	`♧`: [u8(0x83), 0xBD] // U+2667 WHITE CLUB SUIT
	`♣`: [u8(0x83), 0xBE] // U+2663 BLACK CLUB SUIT
	`α`: [u8(0x83), 0xBF] // U+03B1 GREEK SMALL LETTER ALPHA
	`β`: [u8(0x83), 0xC0] // U+03B2 GREEK SMALL LETTER BETA
	`γ`: [u8(0x83), 0xC1] // U+03B3 GREEK SMALL LETTER GAMMA
	`δ`: [u8(0x83), 0xC2] // U+03B4 GREEK SMALL LETTER DELTA
	`ε`: [u8(0x83), 0xC3] // U+03B5 GREEK SMALL LETTER EPSILON
	`ζ`: [u8(0x83), 0xC4] // U+03B6 GREEK SMALL LETTER ZETA
	`η`: [u8(0x83), 0xC5] // U+03B7 GREEK SMALL LETTER ETA
	`θ`: [u8(0x83), 0xC6] // U+03B8 GREEK SMALL LETTER THETA
	`ι`: [u8(0x83), 0xC7] // U+03B9 GREEK SMALL LETTER IOTA
	`κ`: [u8(0x83), 0xC8] // U+03BA GREEK SMALL LETTER KAPPA
	`λ`: [u8(0x83), 0xC9] // U+03BB GREEK SMALL LETTER LAMDA
	`μ`: [u8(0x83), 0xCA] // U+03BC GREEK SMALL LETTER MU
	`ν`: [u8(0x83), 0xCB] // U+03BD GREEK SMALL LETTER NU
	`ξ`: [u8(0x83), 0xCC] // U+03BE GREEK SMALL LETTER XI
	`ο`: [u8(0x83), 0xCD] // U+03BF GREEK SMALL LETTER OMICRON
	`π`: [u8(0x83), 0xCE] // U+03C0 GREEK SMALL LETTER PI
	`ρ`: [u8(0x83), 0xCF] // U+03C1 GREEK SMALL LETTER RHO
	`σ`: [u8(0x83), 0xD0] // U+03C3 GREEK SMALL LETTER SIGMA
	`τ`: [u8(0x83), 0xD1] // U+03C4 GREEK SMALL LETTER TAU
	`υ`: [u8(0x83), 0xD2] // U+03C5 GREEK SMALL LETTER UPSILON
	`φ`: [u8(0x83), 0xD3] // U+03C6 GREEK SMALL LETTER PHI
	`χ`: [u8(0x83), 0xD4] // U+03C7 GREEK SMALL LETTER CHI
	`ψ`: [u8(0x83), 0xD5] // U+03C8 GREEK SMALL LETTER PSI
	`ω`: [u8(0x83), 0xD6] // U+03C9 GREEK SMALL LETTER OMEGA
	`ς`: [u8(0x83), 0xD7] // U+03C2 GREEK SMALL LETTER FINAL SIGMA
	`⓵`: [u8(0x83), 0xD8] // U+24F5 DOUBLE CIRCLED DIGIT ONE
	`⓶`: [u8(0x83), 0xD9] // U+24F6 DOUBLE CIRCLED DIGIT TWO
	`⓷`: [u8(0x83), 0xDA] // U+24F7 DOUBLE CIRCLED DIGIT THREE
	`⓸`: [u8(0x83), 0xDB] // U+24F8 DOUBLE CIRCLED DIGIT FOUR
	`⓹`: [u8(0x83), 0xDC] // U+24F9 DOUBLE CIRCLED DIGIT FIVE
	`⓺`: [u8(0x83), 0xDD] // U+24FA DOUBLE CIRCLED DIGIT SIX
	`⓻`: [u8(0x83), 0xDE] // U+24FB DOUBLE CIRCLED DIGIT SEVEN
	`⓼`: [u8(0x83), 0xDF] // U+24FC DOUBLE CIRCLED DIGIT EIGHT
	`⓽`: [u8(0x83), 0xE0] // U+24FD DOUBLE CIRCLED DIGIT NINE
	`⓾`: [u8(0x83), 0xE1] // U+24FE DOUBLE CIRCLED NUMBER TEN
	`☖`: [u8(0x83), 0xE2] // U+2616 WHITE SHOGI PIECE
	`☗`: [u8(0x83), 0xE3] // U+2617 BLACK SHOGI PIECE
	`〠`: [u8(0x83), 0xE4] // U+3020 POSTAL MARK FACE
	`☎`: [u8(0x83), 0xE5] // U+260E BLACK TELEPHONE
	`☀`: [u8(0x83), 0xE6] // U+2600 BLACK SUN WITH RAYS
	`☁`: [u8(0x83), 0xE7] // U+2601 CLOUD
	`☂`: [u8(0x83), 0xE8] // U+2602 UMBRELLA
	`☃`: [u8(0x83), 0xE9] // U+2603 SNOWMAN
	`♨`: [u8(0x83), 0xEA] // U+2668 HOT SPRINGS
	`▱`: [u8(0x83), 0xEB] // U+25B1 WHITE PARALLELOGRAM
	`ㇰ`: [u8(0x83), 0xEC] // U+31F0 KATAKANA LETTER SMALL KU
	`ㇱ`: [u8(0x83), 0xED] // U+31F1 KATAKANA LETTER SMALL SI
	`ㇲ`: [u8(0x83), 0xEE] // U+31F2 KATAKANA LETTER SMALL SU
	`ㇳ`: [u8(0x83), 0xEF] // U+31F3 KATAKANA LETTER SMALL TO
	`ㇴ`: [u8(0x83), 0xF0] // U+31F4 KATAKANA LETTER SMALL NU
	`ㇵ`: [u8(0x83), 0xF1] // U+31F5 KATAKANA LETTER SMALL HA
	`ㇶ`: [u8(0x83), 0xF2] // U+31F6 KATAKANA LETTER SMALL HI
	`ㇷ`: [u8(0x83), 0xF3] // U+31F7 KATAKANA LETTER SMALL HU
	`ㇸ`: [u8(0x83), 0xF4] // U+31F8 KATAKANA LETTER SMALL HE
	`ㇹ`: [u8(0x83), 0xF5] // U+31F9 KATAKANA LETTER SMALL HO
	`ㇺ`: [u8(0x83), 0xF7] // U+31FA KATAKANA LETTER SMALL MU
	`ㇻ`: [u8(0x83), 0xF8] // U+31FB KATAKANA LETTER SMALL RA
	`ㇼ`: [u8(0x83), 0xF9] // U+31FC KATAKANA LETTER SMALL RI
	`ㇽ`: [u8(0x83), 0xFA] // U+31FD KATAKANA LETTER SMALL RU
	`ㇾ`: [u8(0x83), 0xFB] // U+31FE KATAKANA LETTER SMALL RE
	`ㇿ`: [u8(0x83), 0xFC] // U+31FF KATAKANA LETTER SMALL RO
	`А`: [u8(0x84), 0x40] // U+0410 CYRILLIC CAPITAL LETTER A
	`Б`: [u8(0x84), 0x41] // U+0411 CYRILLIC CAPITAL LETTER BE
	`В`: [u8(0x84), 0x42] // U+0412 CYRILLIC CAPITAL LETTER VE
	`Г`: [u8(0x84), 0x43] // U+0413 CYRILLIC CAPITAL LETTER GHE
	`Д`: [u8(0x84), 0x44] // U+0414 CYRILLIC CAPITAL LETTER DE
	`Е`: [u8(0x84), 0x45] // U+0415 CYRILLIC CAPITAL LETTER IE
	`Ё`: [u8(0x84), 0x46] // U+0401 CYRILLIC CAPITAL LETTER IO
	`Ж`: [u8(0x84), 0x47] // U+0416 CYRILLIC CAPITAL LETTER ZHE
	`З`: [u8(0x84), 0x48] // U+0417 CYRILLIC CAPITAL LETTER ZE
	`И`: [u8(0x84), 0x49] // U+0418 CYRILLIC CAPITAL LETTER I
	`Й`: [u8(0x84), 0x4A] // U+0419 CYRILLIC CAPITAL LETTER SHORT I
	`К`: [u8(0x84), 0x4B] // U+041A CYRILLIC CAPITAL LETTER KA
	`Л`: [u8(0x84), 0x4C] // U+041B CYRILLIC CAPITAL LETTER EL
	`М`: [u8(0x84), 0x4D] // U+041C CYRILLIC CAPITAL LETTER EM
	`Н`: [u8(0x84), 0x4E] // U+041D CYRILLIC CAPITAL LETTER EN
	`О`: [u8(0x84), 0x4F] // U+041E CYRILLIC CAPITAL LETTER O
	`П`: [u8(0x84), 0x50] // U+041F CYRILLIC CAPITAL LETTER PE
	`Р`: [u8(0x84), 0x51] // U+0420 CYRILLIC CAPITAL LETTER ER
	`С`: [u8(0x84), 0x52] // U+0421 CYRILLIC CAPITAL LETTER ES
	`Т`: [u8(0x84), 0x53] // U+0422 CYRILLIC CAPITAL LETTER TE
	`У`: [u8(0x84), 0x54] // U+0423 CYRILLIC CAPITAL LETTER U
	`Ф`: [u8(0x84), 0x55] // U+0424 CYRILLIC CAPITAL LETTER EF
	`Х`: [u8(0x84), 0x56] // U+0425 CYRILLIC CAPITAL LETTER HA
	`Ц`: [u8(0x84), 0x57] // U+0426 CYRILLIC CAPITAL LETTER TSE
	`Ч`: [u8(0x84), 0x58] // U+0427 CYRILLIC CAPITAL LETTER CHE
	`Ш`: [u8(0x84), 0x59] // U+0428 CYRILLIC CAPITAL LETTER SHA
	`Щ`: [u8(0x84), 0x5A] // U+0429 CYRILLIC CAPITAL LETTER SHCHA
	`Ъ`: [u8(0x84), 0x5B] // U+042A CYRILLIC CAPITAL LETTER HARD SIGN
	`Ы`: [u8(0x84), 0x5C] // U+042B CYRILLIC CAPITAL LETTER YERU
	`Ь`: [u8(0x84), 0x5D] // U+042C CYRILLIC CAPITAL LETTER SOFT SIGN
	`Э`: [u8(0x84), 0x5E] // U+042D CYRILLIC CAPITAL LETTER E
	`Ю`: [u8(0x84), 0x5F] // U+042E CYRILLIC CAPITAL LETTER YU
	`Я`: [u8(0x84), 0x60] // U+042F CYRILLIC CAPITAL LETTER YA
	`⎾`: [u8(0x84), 0x61] // U+23BE DENTISTRY SYMBOL LIGHT VERTICAL AND TOP RIGHT
	`⎿`: [u8(0x84), 0x62] // U+23BF DENTISTRY SYMBOL LIGHT VERTICAL AND BOTTOM RIGHT
	`⏀`: [u8(0x84), 0x63] // U+23C0 DENTISTRY SYMBOL LIGHT VERTICAL WITH CIRCLE
	`⏁`: [u8(0x84), 0x64] // U+23C1 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL WITH CIRCLE
	`⏂`: [u8(0x84), 0x65] // U+23C2 DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL WITH CIRCLE
	`⏃`: [u8(0x84), 0x66] // U+23C3 DENTISTRY SYMBOL LIGHT VERTICAL WITH TRIANGLE
	`⏄`: [u8(0x84), 0x67] // U+23C4 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL WITH TRIANGLE
	`⏅`: [u8(0x84), 0x68] // U+23C5 DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL WITH TRIANGLE
	`⏆`: [u8(0x84), 0x69] // U+23C6 DENTISTRY SYMBOL LIGHT VERTICAL AND WAVE
	`⏇`: [u8(0x84), 0x6A] // U+23C7 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL WITH WAVE
	`⏈`: [u8(0x84), 0x6B] // U+23C8 DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL WITH WAVE
	`⏉`: [u8(0x84), 0x6C] // U+23C9 DENTISTRY SYMBOL LIGHT DOWN AND HORIZONTAL
	`⏊`: [u8(0x84), 0x6D] // U+23CA DENTISTRY SYMBOL LIGHT UP AND HORIZONTAL
	`⏋`: [u8(0x84), 0x6E] // U+23CB DENTISTRY SYMBOL LIGHT VERTICAL AND TOP LEFT
	`⏌`: [u8(0x84), 0x6F] // U+23CC DENTISTRY SYMBOL LIGHT VERTICAL AND BOTTOM LEFT
	`а`: [u8(0x84), 0x70] // U+0430 CYRILLIC SMALL LETTER A
	`б`: [u8(0x84), 0x71] // U+0431 CYRILLIC SMALL LETTER BE
	`в`: [u8(0x84), 0x72] // U+0432 CYRILLIC SMALL LETTER VE
	`г`: [u8(0x84), 0x73] // U+0433 CYRILLIC SMALL LETTER GHE
	`д`: [u8(0x84), 0x74] // U+0434 CYRILLIC SMALL LETTER DE
	`е`: [u8(0x84), 0x75] // U+0435 CYRILLIC SMALL LETTER IE
	`ё`: [u8(0x84), 0x76] // U+0451 CYRILLIC SMALL LETTER IO
	`ж`: [u8(0x84), 0x77] // U+0436 CYRILLIC SMALL LETTER ZHE
	`з`: [u8(0x84), 0x78] // U+0437 CYRILLIC SMALL LETTER ZE
	`и`: [u8(0x84), 0x79] // U+0438 CYRILLIC SMALL LETTER I
	`й`: [u8(0x84), 0x7A] // U+0439 CYRILLIC SMALL LETTER SHORT I
	`к`: [u8(0x84), 0x7B] // U+043A CYRILLIC SMALL LETTER KA
	`л`: [u8(0x84), 0x7C] // U+043B CYRILLIC SMALL LETTER EL
	`м`: [u8(0x84), 0x7D] // U+043C CYRILLIC SMALL LETTER EM
	`н`: [u8(0x84), 0x7E] // U+043D CYRILLIC SMALL LETTER EN
	`о`: [u8(0x84), 0x80] // U+043E CYRILLIC SMALL LETTER O
	`п`: [u8(0x84), 0x81] // U+043F CYRILLIC SMALL LETTER PE
	`р`: [u8(0x84), 0x82] // U+0440 CYRILLIC SMALL LETTER ER
	`с`: [u8(0x84), 0x83] // U+0441 CYRILLIC SMALL LETTER ES
	`т`: [u8(0x84), 0x84] // U+0442 CYRILLIC SMALL LETTER TE
	`у`: [u8(0x84), 0x85] // U+0443 CYRILLIC SMALL LETTER U
	`ф`: [u8(0x84), 0x86] // U+0444 CYRILLIC SMALL LETTER EF
	`х`: [u8(0x84), 0x87] // U+0445 CYRILLIC SMALL LETTER HA
	`ц`: [u8(0x84), 0x88] // U+0446 CYRILLIC SMALL LETTER TSE
	`ч`: [u8(0x84), 0x89] // U+0447 CYRILLIC SMALL LETTER CHE
	`ш`: [u8(0x84), 0x8A] // U+0448 CYRILLIC SMALL LETTER SHA
	`щ`: [u8(0x84), 0x8B] // U+0449 CYRILLIC SMALL LETTER SHCHA
	`ъ`: [u8(0x84), 0x8C] // U+044A CYRILLIC SMALL LETTER HARD SIGN
	`ы`: [u8(0x84), 0x8D] // U+044B CYRILLIC SMALL LETTER YERU
	`ь`: [u8(0x84), 0x8E] // U+044C CYRILLIC SMALL LETTER SOFT SIGN
	`э`: [u8(0x84), 0x8F] // U+044D CYRILLIC SMALL LETTER E
	`ю`: [u8(0x84), 0x90] // U+044E CYRILLIC SMALL LETTER YU
	`я`: [u8(0x84), 0x91] // U+044F CYRILLIC SMALL LETTER YA
	`ヷ`: [u8(0x84), 0x92] // U+30F7 KATAKANA LETTER VA
	`ヸ`: [u8(0x84), 0x93] // U+30F8 KATAKANA LETTER VI
	`ヹ`: [u8(0x84), 0x94] // U+30F9 KATAKANA LETTER VE
	`ヺ`: [u8(0x84), 0x95] // U+30FA KATAKANA LETTER VO
	`⋚`: [u8(0x84), 0x96] // U+22DA LESS-THAN EQUAL TO OR GREATER-THAN
	`⋛`: [u8(0x84), 0x97] // U+22DB GREATER-THAN EQUAL TO OR LESS-THAN
	`⅓`: [u8(0x84), 0x98] // U+2153 VULGAR FRACTION ONE THIRD
	`⅔`: [u8(0x84), 0x99] // U+2154 VULGAR FRACTION TWO THIRDS
	`⅕`: [u8(0x84), 0x9A] // U+2155 VULGAR FRACTION ONE FIFTH
	`✓`: [u8(0x84), 0x9B] // U+2713 CHECK MARK
	`⌘`: [u8(0x84), 0x9C] // U+2318 PLACE OF INTEREST SIGN
	`␣`: [u8(0x84), 0x9D] // U+2423 OPEN BOX
	`⏎`: [u8(0x84), 0x9E] // U+23CE RETURN SYMBOL
	`─`: [u8(0x84), 0x9F] // U+2500 BOX DRAWINGS LIGHT HORIZONTAL
	`│`: [u8(0x84), 0xA0] // U+2502 BOX DRAWINGS LIGHT VERTICAL
	`┌`: [u8(0x84), 0xA1] // U+250C BOX DRAWINGS LIGHT DOWN AND RIGHT
	`┐`: [u8(0x84), 0xA2] // U+2510 BOX DRAWINGS LIGHT DOWN AND LEFT
	`┘`: [u8(0x84), 0xA3] // U+2518 BOX DRAWINGS LIGHT UP AND LEFT
	`└`: [u8(0x84), 0xA4] // U+2514 BOX DRAWINGS LIGHT UP AND RIGHT
	`├`: [u8(0x84), 0xA5] // U+251C BOX DRAWINGS LIGHT VERTICAL AND RIGHT
	`┬`: [u8(0x84), 0xA6] // U+252C BOX DRAWINGS LIGHT DOWN AND HORIZONTAL
	`┤`: [u8(0x84), 0xA7] // U+2524 BOX DRAWINGS LIGHT VERTICAL AND LEFT
	`┴`: [u8(0x84), 0xA8] // U+2534 BOX DRAWINGS LIGHT UP AND HORIZONTAL
	`┼`: [u8(0x84), 0xA9] // U+253C BOX DRAWINGS LIGHT VERTICAL AND HORIZONTAL
	`━`: [u8(0x84), 0xAA] // U+2501 BOX DRAWINGS HEAVY HORIZONTAL
	`┃`: [u8(0x84), 0xAB] // U+2503 BOX DRAWINGS HEAVY VERTICAL
	`┏`: [u8(0x84), 0xAC] // U+250F BOX DRAWINGS HEAVY DOWN AND RIGHT
	`┓`: [u8(0x84), 0xAD] // U+2513 BOX DRAWINGS HEAVY DOWN AND LEFT
	`┛`: [u8(0x84), 0xAE] // U+251B BOX DRAWINGS HEAVY UP AND LEFT
	`┗`: [u8(0x84), 0xAF] // U+2517 BOX DRAWINGS HEAVY UP AND RIGHT
	`┣`: [u8(0x84), 0xB0] // U+2523 BOX DRAWINGS HEAVY VERTICAL AND RIGHT
	`┳`: [u8(0x84), 0xB1] // U+2533 BOX DRAWINGS HEAVY DOWN AND HORIZONTAL
	`┫`: [u8(0x84), 0xB2] // U+252B BOX DRAWINGS HEAVY VERTICAL AND LEFT
	`┻`: [u8(0x84), 0xB3] // U+253B BOX DRAWINGS HEAVY UP AND HORIZONTAL
	`╋`: [u8(0x84), 0xB4] // U+254B BOX DRAWINGS HEAVY VERTICAL AND HORIZONTAL
	`┠`: [u8(0x84), 0xB5] // U+2520 BOX DRAWINGS VERTICAL HEAVY AND RIGHT LIGHT
	`┯`: [u8(0x84), 0xB6] // U+252F BOX DRAWINGS DOWN LIGHT AND HORIZONTAL HEAVY
	`┨`: [u8(0x84), 0xB7] // U+2528 BOX DRAWINGS VERTICAL HEAVY AND LEFT LIGHT
	`┷`: [u8(0x84), 0xB8] // U+2537 BOX DRAWINGS UP LIGHT AND HORIZONTAL HEAVY
	`┿`: [u8(0x84), 0xB9] // U+253F BOX DRAWINGS VERTICAL LIGHT AND HORIZONTAL HEAVY
	`┝`: [u8(0x84), 0xBA] // U+251D BOX DRAWINGS VERTICAL LIGHT AND RIGHT HEAVY
	`┰`: [u8(0x84), 0xBB] // U+2530 BOX DRAWINGS DOWN HEAVY AND HORIZONTAL LIGHT
	`┥`: [u8(0x84), 0xBC] // U+2525 BOX DRAWINGS VERTICAL LIGHT AND LEFT HEAVY
	`┸`: [u8(0x84), 0xBD] // U+2538 BOX DRAWINGS UP HEAVY AND HORIZONTAL LIGHT
	`╂`: [u8(0x84), 0xBE] // U+2542 BOX DRAWINGS VERTICAL HEAVY AND HORIZONTAL LIGHT
	`㉑`: [u8(0x84), 0xBF] // U+3251 CIRCLED NUMBER TWENTY ONE
	`㉒`: [u8(0x84), 0xC0] // U+3252 CIRCLED NUMBER TWENTY TWO
	`㉓`: [u8(0x84), 0xC1] // U+3253 CIRCLED NUMBER TWENTY THREE
	`㉔`: [u8(0x84), 0xC2] // U+3254 CIRCLED NUMBER TWENTY FOUR
	`㉕`: [u8(0x84), 0xC3] // U+3255 CIRCLED NUMBER TWENTY FIVE
	`㉖`: [u8(0x84), 0xC4] // U+3256 CIRCLED NUMBER TWENTY SIX
	`㉗`: [u8(0x84), 0xC5] // U+3257 CIRCLED NUMBER TWENTY SEVEN
	`㉘`: [u8(0x84), 0xC6] // U+3258 CIRCLED NUMBER TWENTY EIGHT
	`㉙`: [u8(0x84), 0xC7] // U+3259 CIRCLED NUMBER TWENTY NINE
	`㉚`: [u8(0x84), 0xC8] // U+325A CIRCLED NUMBER THIRTY
	`㉛`: [u8(0x84), 0xC9] // U+325B CIRCLED NUMBER THIRTY ONE
	`㉜`: [u8(0x84), 0xCA] // U+325C CIRCLED NUMBER THIRTY TWO
	`㉝`: [u8(0x84), 0xCB] // U+325D CIRCLED NUMBER THIRTY THREE
	`㉞`: [u8(0x84), 0xCC] // U+325E CIRCLED NUMBER THIRTY FOUR
	`㉟`: [u8(0x84), 0xCD] // U+325F CIRCLED NUMBER THIRTY FIVE
	`㊱`: [u8(0x84), 0xCE] // U+32B1 CIRCLED NUMBER THIRTY SIX
	`㊲`: [u8(0x84), 0xCF] // U+32B2 CIRCLED NUMBER THIRTY SEVEN
	`㊳`: [u8(0x84), 0xD0] // U+32B3 CIRCLED NUMBER THIRTY EIGHT
	`㊴`: [u8(0x84), 0xD1] // U+32B4 CIRCLED NUMBER THIRTY NINE
	`㊵`: [u8(0x84), 0xD2] // U+32B5 CIRCLED NUMBER FORTY
	`㊶`: [u8(0x84), 0xD3] // U+32B6 CIRCLED NUMBER FORTY ONE
	`㊷`: [u8(0x84), 0xD4] // U+32B7 CIRCLED NUMBER FORTY TWO
	`㊸`: [u8(0x84), 0xD5] // U+32B8 CIRCLED NUMBER FORTY THREE
	`㊹`: [u8(0x84), 0xD6] // U+32B9 CIRCLED NUMBER FORTY FOUR
	`㊺`: [u8(0x84), 0xD7] // U+32BA CIRCLED NUMBER FORTY FIVE
	`㊻`: [u8(0x84), 0xD8] // U+32BB CIRCLED NUMBER FORTY SIX
	`㊼`: [u8(0x84), 0xD9] // U+32BC CIRCLED NUMBER FORTY SEVEN
	`㊽`: [u8(0x84), 0xDA] // U+32BD CIRCLED NUMBER FORTY EIGHT
	`㊾`: [u8(0x84), 0xDB] // U+32BE CIRCLED NUMBER FORTY NINE
	`㊿`: [u8(0x84), 0xDC] // U+32BF CIRCLED NUMBER FIFTY
	`◐`: [u8(0x84), 0xE5] // U+25D0 CIRCLE WITH LEFT HALF BLACK
	`◑`: [u8(0x84), 0xE6] // U+25D1 CIRCLE WITH RIGHT HALF BLACK
	`◒`: [u8(0x84), 0xE7] // U+25D2 CIRCLE WITH LOWER HALF BLACK
	`◓`: [u8(0x84), 0xE8] // U+25D3 CIRCLE WITH UPPER HALF BLACK
	`‼`: [u8(0x84), 0xE9] // U+203C DOUBLE EXCLAMATION MARK
	`⁇`: [u8(0x84), 0xEA] // U+2047 DOUBLE QUESTION MARK
	`⁈`: [u8(0x84), 0xEB] // U+2048 QUESTION EXCLAMATION MARK
	`⁉`: [u8(0x84), 0xEC] // U+2049 EXCLAMATION QUESTION MARK
	`Ǎ`: [u8(0x84), 0xED] // U+01CD LATIN CAPITAL LETTER A WITH CARON
	`ǎ`: [u8(0x84), 0xEE] // U+01CE LATIN SMALL LETTER A WITH CARON
	`ǐ`: [u8(0x84), 0xEF] // U+01D0 LATIN SMALL LETTER I WITH CARON
	`Ḿ`: [u8(0x84), 0xF0] // U+1E3E LATIN CAPITAL LETTER M WITH ACUTE
	`ḿ`: [u8(0x84), 0xF1] // U+1E3F LATIN SMALL LETTER M WITH ACUTE
	`Ǹ`: [u8(0x84), 0xF2] // U+01F8 LATIN CAPITAL LETTER N WITH GRAVE
	`ǹ`: [u8(0x84), 0xF3] // U+01F9 LATIN SMALL LETTER N WITH GRAVE
	`Ǒ`: [u8(0x84), 0xF4] // U+01D1 LATIN CAPITAL LETTER O WITH CARON
	`ǒ`: [u8(0x84), 0xF5] // U+01D2 LATIN SMALL LETTER O WITH CARON
	`ǔ`: [u8(0x84), 0xF6] // U+01D4 LATIN SMALL LETTER U WITH CARON
	`ǖ`: [u8(0x84), 0xF7] // U+01D6 LATIN SMALL LETTER U WITH DIAERESIS AND MACRON
	`ǘ`: [u8(0x84), 0xF8] // U+01D8 LATIN SMALL LETTER U WITH DIAERESIS AND ACUTE
	`ǚ`: [u8(0x84), 0xF9] // U+01DA LATIN SMALL LETTER U WITH DIAERESIS AND CARON
	`ǜ`: [u8(0x84), 0xFA] // U+01DC LATIN SMALL LETTER U WITH DIAERESIS AND GRAVE
	`€`: [u8(0x85), 0x40] // U+20AC EURO SIGN
	` `: [u8(0x85), 0x41] // U+00A0 NO-BREAK SPACE
	`¡`: [u8(0x85), 0x42] // U+00A1 INVERTED EXCLAMATION MARK
	`¤`: [u8(0x85), 0x43] // U+00A4 CURRENCY SIGN
	`¦`: [u8(0x85), 0x44] // U+00A6 BROKEN BAR
	`©`: [u8(0x85), 0x45] // U+00A9 COPYRIGHT SIGN
	`ª`: [u8(0x85), 0x46] // U+00AA FEMININE ORDINAL INDICATOR
	`«`: [u8(0x85), 0x47] // U+00AB LEFT-POINTING DOUBLE ANGLE QUOTATION MARK
	`­`: [u8(0x85), 0x48] // U+00AD SOFT HYPHEN
	`®`: [u8(0x85), 0x49] // U+00AE REGISTERED SIGN
	`¯`: [u8(0x85), 0x4A] // U+00AF MACRON
	`²`: [u8(0x85), 0x4B] // U+00B2 SUPERSCRIPT TWO
	`³`: [u8(0x85), 0x4C] // U+00B3 SUPERSCRIPT THREE
	`·`: [u8(0x85), 0x4D] // U+00B7 MIDDLE DOT
	`¸`: [u8(0x85), 0x4E] // U+00B8 CEDILLA
	`¹`: [u8(0x85), 0x4F] // U+00B9 SUPERSCRIPT ONE
	`º`: [u8(0x85), 0x50] // U+00BA MASCULINE ORDINAL INDICATOR
	`»`: [u8(0x85), 0x51] // U+00BB RIGHT-POINTING DOUBLE ANGLE QUOTATION MARK
	`¼`: [u8(0x85), 0x52] // U+00BC VULGAR FRACTION ONE QUARTER
	`½`: [u8(0x85), 0x53] // U+00BD VULGAR FRACTION ONE HALF
	`¾`: [u8(0x85), 0x54] // U+00BE VULGAR FRACTION THREE QUARTERS
	`¿`: [u8(0x85), 0x55] // U+00BF INVERTED QUESTION MARK
	`À`: [u8(0x85), 0x56] // U+00C0 LATIN CAPITAL LETTER A WITH GRAVE
	`Á`: [u8(0x85), 0x57] // U+00C1 LATIN CAPITAL LETTER A WITH ACUTE
	`Â`: [u8(0x85), 0x58] // U+00C2 LATIN CAPITAL LETTER A WITH CIRCUMFLEX
	`Ã`: [u8(0x85), 0x59] // U+00C3 LATIN CAPITAL LETTER A WITH TILDE
	`Ä`: [u8(0x85), 0x5A] // U+00C4 LATIN CAPITAL LETTER A WITH DIAERESIS
	`Å`: [u8(0x85), 0x5B] // U+00C5 LATIN CAPITAL LETTER A WITH RING ABOVE
	`Æ`: [u8(0x85), 0x5C] // U+00C6 LATIN CAPITAL LETTER AE
	`Ç`: [u8(0x85), 0x5D] // U+00C7 LATIN CAPITAL LETTER C WITH CEDILLA
	`È`: [u8(0x85), 0x5E] // U+00C8 LATIN CAPITAL LETTER E WITH GRAVE
	`É`: [u8(0x85), 0x5F] // U+00C9 LATIN CAPITAL LETTER E WITH ACUTE
	`Ê`: [u8(0x85), 0x60] // U+00CA LATIN CAPITAL LETTER E WITH CIRCUMFLEX
	`Ë`: [u8(0x85), 0x61] // U+00CB LATIN CAPITAL LETTER E WITH DIAERESIS
	`Ì`: [u8(0x85), 0x62] // U+00CC LATIN CAPITAL LETTER I WITH GRAVE
	`Í`: [u8(0x85), 0x63] // U+00CD LATIN CAPITAL LETTER I WITH ACUTE
	`Î`: [u8(0x85), 0x64] // U+00CE LATIN CAPITAL LETTER I WITH CIRCUMFLEX
	`Ï`: [u8(0x85), 0x65] // U+00CF LATIN CAPITAL LETTER I WITH DIAERESIS
	`Ð`: [u8(0x85), 0x66] // U+00D0 LATIN CAPITAL LETTER ETH
	`Ñ`: [u8(0x85), 0x67] // U+00D1 LATIN CAPITAL LETTER N WITH TILDE
	`Ò`: [u8(0x85), 0x68] // U+00D2 LATIN CAPITAL LETTER O WITH GRAVE
	`Ó`: [u8(0x85), 0x69] // U+00D3 LATIN CAPITAL LETTER O WITH ACUTE
	`Ô`: [u8(0x85), 0x6A] // U+00D4 LATIN CAPITAL LETTER O WITH CIRCUMFLEX
	`Õ`: [u8(0x85), 0x6B] // U+00D5 LATIN CAPITAL LETTER O WITH TILDE
	`Ö`: [u8(0x85), 0x6C] // U+00D6 LATIN CAPITAL LETTER O WITH DIAERESIS
	`Ø`: [u8(0x85), 0x6D] // U+00D8 LATIN CAPITAL LETTER O WITH STROKE
	`Ù`: [u8(0x85), 0x6E] // U+00D9 LATIN CAPITAL LETTER U WITH GRAVE
	`Ú`: [u8(0x85), 0x6F] // U+00DA LATIN CAPITAL LETTER U WITH ACUTE
	`Û`: [u8(0x85), 0x70] // U+00DB LATIN CAPITAL LETTER U WITH CIRCUMFLEX
	`Ü`: [u8(0x85), 0x71] // U+00DC LATIN CAPITAL LETTER U WITH DIAERESIS
	`Ý`: [u8(0x85), 0x72] // U+00DD LATIN CAPITAL LETTER Y WITH ACUTE
	`Þ`: [u8(0x85), 0x73] // U+00DE LATIN CAPITAL LETTER THORN
	`ß`: [u8(0x85), 0x74] // U+00DF LATIN SMALL LETTER SHARP S
	`à`: [u8(0x85), 0x75] // U+00E0 LATIN SMALL LETTER A WITH GRAVE
	`á`: [u8(0x85), 0x76] // U+00E1 LATIN SMALL LETTER A WITH ACUTE
	`â`: [u8(0x85), 0x77] // U+00E2 LATIN SMALL LETTER A WITH CIRCUMFLEX
	`ã`: [u8(0x85), 0x78] // U+00E3 LATIN SMALL LETTER A WITH TILDE
	`ä`: [u8(0x85), 0x79] // U+00E4 LATIN SMALL LETTER A WITH DIAERESIS
	`å`: [u8(0x85), 0x7A] // U+00E5 LATIN SMALL LETTER A WITH RING ABOVE
	`æ`: [u8(0x85), 0x7B] // U+00E6 LATIN SMALL LETTER AE
	`ç`: [u8(0x85), 0x7C] // U+00E7 LATIN SMALL LETTER C WITH CEDILLA
	`è`: [u8(0x85), 0x7D] // U+00E8 LATIN SMALL LETTER E WITH GRAVE
	`é`: [u8(0x85), 0x7E] // U+00E9 LATIN SMALL LETTER E WITH ACUTE
	`ê`: [u8(0x85), 0x80] // U+00EA LATIN SMALL LETTER E WITH CIRCUMFLEX
	`ë`: [u8(0x85), 0x81] // U+00EB LATIN SMALL LETTER E WITH DIAERESIS
	`ì`: [u8(0x85), 0x82] // U+00EC LATIN SMALL LETTER I WITH GRAVE
	`í`: [u8(0x85), 0x83] // U+00ED LATIN SMALL LETTER I WITH ACUTE
	`î`: [u8(0x85), 0x84] // U+00EE LATIN SMALL LETTER I WITH CIRCUMFLEX
	`ï`: [u8(0x85), 0x85] // U+00EF LATIN SMALL LETTER I WITH DIAERESIS
	`ð`: [u8(0x85), 0x86] // U+00F0 LATIN SMALL LETTER ETH
	`ñ`: [u8(0x85), 0x87] // U+00F1 LATIN SMALL LETTER N WITH TILDE
	`ò`: [u8(0x85), 0x88] // U+00F2 LATIN SMALL LETTER O WITH GRAVE
	`ó`: [u8(0x85), 0x89] // U+00F3 LATIN SMALL LETTER O WITH ACUTE
	`ô`: [u8(0x85), 0x8A] // U+00F4 LATIN SMALL LETTER O WITH CIRCUMFLEX
	`õ`: [u8(0x85), 0x8B] // U+00F5 LATIN SMALL LETTER O WITH TILDE
	`ö`: [u8(0x85), 0x8C] // U+00F6 LATIN SMALL LETTER O WITH DIAERESIS
	`ø`: [u8(0x85), 0x8D] // U+00F8 LATIN SMALL LETTER O WITH STROKE
	`ù`: [u8(0x85), 0x8E] // U+00F9 LATIN SMALL LETTER U WITH GRAVE
	`ú`: [u8(0x85), 0x8F] // U+00FA LATIN SMALL LETTER U WITH ACUTE
	`û`: [u8(0x85), 0x90] // U+00FB LATIN SMALL LETTER U WITH CIRCUMFLEX
	`ü`: [u8(0x85), 0x91] // U+00FC LATIN SMALL LETTER U WITH DIAERESIS
	`ý`: [u8(0x85), 0x92] // U+00FD LATIN SMALL LETTER Y WITH ACUTE
	`þ`: [u8(0x85), 0x93] // U+00FE LATIN SMALL LETTER THORN
	`ÿ`: [u8(0x85), 0x94] // U+00FF LATIN SMALL LETTER Y WITH DIAERESIS
	`Ā`: [u8(0x85), 0x95] // U+0100 LATIN CAPITAL LETTER A WITH MACRON
	`Ī`: [u8(0x85), 0x96] // U+012A LATIN CAPITAL LETTER I WITH MACRON
	`Ū`: [u8(0x85), 0x97] // U+016A LATIN CAPITAL LETTER U WITH MACRON
	`Ē`: [u8(0x85), 0x98] // U+0112 LATIN CAPITAL LETTER E WITH MACRON
	`Ō`: [u8(0x85), 0x99] // U+014C LATIN CAPITAL LETTER O WITH MACRON
	`ā`: [u8(0x85), 0x9A] // U+0101 LATIN SMALL LETTER A WITH MACRON
	`ī`: [u8(0x85), 0x9B] // U+012B LATIN SMALL LETTER I WITH MACRON
	`ū`: [u8(0x85), 0x9C] // U+016B LATIN SMALL LETTER U WITH MACRON
	`ē`: [u8(0x85), 0x9D] // U+0113 LATIN SMALL LETTER E WITH MACRON
	`ō`: [u8(0x85), 0x9E] // U+014D LATIN SMALL LETTER O WITH MACRON
	`Ą`: [u8(0x85), 0x9F] // U+0104 LATIN CAPITAL LETTER A WITH OGONEK
	`˘`: [u8(0x85), 0xA0] // U+02D8 BREVE
	`Ł`: [u8(0x85), 0xA1] // U+0141 LATIN CAPITAL LETTER L WITH STROKE
	`Ľ`: [u8(0x85), 0xA2] // U+013D LATIN CAPITAL LETTER L WITH CARON
	`Ś`: [u8(0x85), 0xA3] // U+015A LATIN CAPITAL LETTER S WITH ACUTE
	`Š`: [u8(0x85), 0xA4] // U+0160 LATIN CAPITAL LETTER S WITH CARON
	`Ş`: [u8(0x85), 0xA5] // U+015E LATIN CAPITAL LETTER S WITH CEDILLA
	`Ť`: [u8(0x85), 0xA6] // U+0164 LATIN CAPITAL LETTER T WITH CARON
	`Ź`: [u8(0x85), 0xA7] // U+0179 LATIN CAPITAL LETTER Z WITH ACUTE
	`Ž`: [u8(0x85), 0xA8] // U+017D LATIN CAPITAL LETTER Z WITH CARON
	`Ż`: [u8(0x85), 0xA9] // U+017B LATIN CAPITAL LETTER Z WITH DOT ABOVE
	`ą`: [u8(0x85), 0xAA] // U+0105 LATIN SMALL LETTER A WITH OGONEK
	`˛`: [u8(0x85), 0xAB] // U+02DB OGONEK
	`ł`: [u8(0x85), 0xAC] // U+0142 LATIN SMALL LETTER L WITH STROKE
	`ľ`: [u8(0x85), 0xAD] // U+013E LATIN SMALL LETTER L WITH CARON
	`ś`: [u8(0x85), 0xAE] // U+015B LATIN SMALL LETTER S WITH ACUTE
	`ˇ`: [u8(0x85), 0xAF] // U+02C7 CARON
	`š`: [u8(0x85), 0xB0] // U+0161 LATIN SMALL LETTER S WITH CARON
	`ş`: [u8(0x85), 0xB1] // U+015F LATIN SMALL LETTER S WITH CEDILLA
	`ť`: [u8(0x85), 0xB2] // U+0165 LATIN SMALL LETTER T WITH CARON
	`ź`: [u8(0x85), 0xB3] // U+017A LATIN SMALL LETTER Z WITH ACUTE
	`˝`: [u8(0x85), 0xB4] // U+02DD DOUBLE ACUTE ACCENT
	`ž`: [u8(0x85), 0xB5] // U+017E LATIN SMALL LETTER Z WITH CARON
	`ż`: [u8(0x85), 0xB6] // U+017C LATIN SMALL LETTER Z WITH DOT ABOVE
	`Ŕ`: [u8(0x85), 0xB7] // U+0154 LATIN CAPITAL LETTER R WITH ACUTE
	`Ă`: [u8(0x85), 0xB8] // U+0102 LATIN CAPITAL LETTER A WITH BREVE
	`Ĺ`: [u8(0x85), 0xB9] // U+0139 LATIN CAPITAL LETTER L WITH ACUTE
	`Ć`: [u8(0x85), 0xBA] // U+0106 LATIN CAPITAL LETTER C WITH ACUTE
	`Č`: [u8(0x85), 0xBB] // U+010C LATIN CAPITAL LETTER C WITH CARON
	`Ę`: [u8(0x85), 0xBC] // U+0118 LATIN CAPITAL LETTER E WITH OGONEK
	`Ě`: [u8(0x85), 0xBD] // U+011A LATIN CAPITAL LETTER E WITH CARON
	`Ď`: [u8(0x85), 0xBE] // U+010E LATIN CAPITAL LETTER D WITH CARON
	`Ń`: [u8(0x85), 0xBF] // U+0143 LATIN CAPITAL LETTER N WITH ACUTE
	`Ň`: [u8(0x85), 0xC0] // U+0147 LATIN CAPITAL LETTER N WITH CARON
	`Ő`: [u8(0x85), 0xC1] // U+0150 LATIN CAPITAL LETTER O WITH DOUBLE ACUTE
	`Ř`: [u8(0x85), 0xC2] // U+0158 LATIN CAPITAL LETTER R WITH CARON
	`Ů`: [u8(0x85), 0xC3] // U+016E LATIN CAPITAL LETTER U WITH RING ABOVE
	`Ű`: [u8(0x85), 0xC4] // U+0170 LATIN CAPITAL LETTER U WITH DOUBLE ACUTE
	`Ţ`: [u8(0x85), 0xC5] // U+0162 LATIN CAPITAL LETTER T WITH CEDILLA
	`ŕ`: [u8(0x85), 0xC6] // U+0155 LATIN SMALL LETTER R WITH ACUTE
	`ă`: [u8(0x85), 0xC7] // U+0103 LATIN SMALL LETTER A WITH BREVE
	`ĺ`: [u8(0x85), 0xC8] // U+013A LATIN SMALL LETTER L WITH ACUTE
	`ć`: [u8(0x85), 0xC9] // U+0107 LATIN SMALL LETTER C WITH ACUTE
	`č`: [u8(0x85), 0xCA] // U+010D LATIN SMALL LETTER C WITH CARON
	`ę`: [u8(0x85), 0xCB] // U+0119 LATIN SMALL LETTER E WITH OGONEK
	`ě`: [u8(0x85), 0xCC] // U+011B LATIN SMALL LETTER E WITH CARON
	`ď`: [u8(0x85), 0xCD] // U+010F LATIN SMALL LETTER D WITH CARON
	`đ`: [u8(0x85), 0xCE] // U+0111 LATIN SMALL LETTER D WITH STROKE
	`ń`: [u8(0x85), 0xCF] // U+0144 LATIN SMALL LETTER N WITH ACUTE
	`ň`: [u8(0x85), 0xD0] // U+0148 LATIN SMALL LETTER N WITH CARON
	`ő`: [u8(0x85), 0xD1] // U+0151 LATIN SMALL LETTER O WITH DOUBLE ACUTE
	`ř`: [u8(0x85), 0xD2] // U+0159 LATIN SMALL LETTER R WITH CARON
	`ů`: [u8(0x85), 0xD3] // U+016F LATIN SMALL LETTER U WITH RING ABOVE
	`ű`: [u8(0x85), 0xD4] // U+0171 LATIN SMALL LETTER U WITH DOUBLE ACUTE
	`ţ`: [u8(0x85), 0xD5] // U+0163 LATIN SMALL LETTER T WITH CEDILLA
	`˙`: [u8(0x85), 0xD6] // U+02D9 DOT ABOVE
	`Ĉ`: [u8(0x85), 0xD7] // U+0108 LATIN CAPITAL LETTER C WITH CIRCUMFLEX
	`Ĝ`: [u8(0x85), 0xD8] // U+011C LATIN CAPITAL LETTER G WITH CIRCUMFLEX
	`Ĥ`: [u8(0x85), 0xD9] // U+0124 LATIN CAPITAL LETTER H WITH CIRCUMFLEX
	`Ĵ`: [u8(0x85), 0xDA] // U+0134 LATIN CAPITAL LETTER J WITH CIRCUMFLEX
	`Ŝ`: [u8(0x85), 0xDB] // U+015C LATIN CAPITAL LETTER S WITH CIRCUMFLEX
	`Ŭ`: [u8(0x85), 0xDC] // U+016C LATIN CAPITAL LETTER U WITH BREVE
	`ĉ`: [u8(0x85), 0xDD] // U+0109 LATIN SMALL LETTER C WITH CIRCUMFLEX
	`ĝ`: [u8(0x85), 0xDE] // U+011D LATIN SMALL LETTER G WITH CIRCUMFLEX
	`ĥ`: [u8(0x85), 0xDF] // U+0125 LATIN SMALL LETTER H WITH CIRCUMFLEX
	`ĵ`: [u8(0x85), 0xE0] // U+0135 LATIN SMALL LETTER J WITH CIRCUMFLEX
	`ŝ`: [u8(0x85), 0xE1] // U+015D LATIN SMALL LETTER S WITH CIRCUMFLEX
	`ŭ`: [u8(0x85), 0xE2] // U+016D LATIN SMALL LETTER U WITH BREVE
	`ɱ`: [u8(0x85), 0xE3] // U+0271 LATIN SMALL LETTER M WITH HOOK
	`ʋ`: [u8(0x85), 0xE4] // U+028B LATIN SMALL LETTER V WITH HOOK
	`ɾ`: [u8(0x85), 0xE5] // U+027E LATIN SMALL LETTER R WITH FISHHOOK
	`ʃ`: [u8(0x85), 0xE6] // U+0283 LATIN SMALL LETTER ESH
	`ʒ`: [u8(0x85), 0xE7] // U+0292 LATIN SMALL LETTER EZH
	`ɬ`: [u8(0x85), 0xE8] // U+026C LATIN SMALL LETTER L WITH BELT
	`ɮ`: [u8(0x85), 0xE9] // U+026E LATIN SMALL LETTER LEZH
	`ɹ`: [u8(0x85), 0xEA] // U+0279 LATIN SMALL LETTER TURNED R
	`ʈ`: [u8(0x85), 0xEB] // U+0288 LATIN SMALL LETTER T WITH RETROFLEX HOOK
	`ɖ`: [u8(0x85), 0xEC] // U+0256 LATIN SMALL LETTER D WITH TAIL
	`ɳ`: [u8(0x85), 0xED] // U+0273 LATIN SMALL LETTER N WITH RETROFLEX HOOK
	`ɽ`: [u8(0x85), 0xEE] // U+027D LATIN SMALL LETTER R WITH TAIL
	`ʂ`: [u8(0x85), 0xEF] // U+0282 LATIN SMALL LETTER S WITH HOOK
	`ʐ`: [u8(0x85), 0xF0] // U+0290 LATIN SMALL LETTER Z WITH RETROFLEX HOOK
	`ɻ`: [u8(0x85), 0xF1] // U+027B LATIN SMALL LETTER TURNED R WITH HOOK
	`ɭ`: [u8(0x85), 0xF2] // U+026D LATIN SMALL LETTER L WITH RETROFLEX HOOK
	`ɟ`: [u8(0x85), 0xF3] // U+025F LATIN SMALL LETTER DOTLESS J WITH STROKE
	`ɲ`: [u8(0x85), 0xF4] // U+0272 LATIN SMALL LETTER N WITH LEFT HOOK
	`ʝ`: [u8(0x85), 0xF5] // U+029D LATIN SMALL LETTER J WITH CROSSED-TAIL
	`ʎ`: [u8(0x85), 0xF6] // U+028E LATIN SMALL LETTER TURNED Y
	`ɡ`: [u8(0x85), 0xF7] // U+0261 LATIN SMALL LETTER SCRIPT G
	`ŋ`: [u8(0x85), 0xF8] // U+014B LATIN SMALL LETTER ENG
	`ɰ`: [u8(0x85), 0xF9] // U+0270 LATIN SMALL LETTER TURNED M WITH LONG LEG
	`ʁ`: [u8(0x85), 0xFA] // U+0281 LATIN LETTER SMALL CAPITAL INVERTED R
	`ħ`: [u8(0x85), 0xFB] // U+0127 LATIN SMALL LETTER H WITH STROKE
	`ʕ`: [u8(0x85), 0xFC] // U+0295 LATIN LETTER PHARYNGEAL VOICED FRICATIVE
	`ʔ`: [u8(0x86), 0x40] // U+0294 LATIN LETTER GLOTTAL STOP
	`ɦ`: [u8(0x86), 0x41] // U+0266 LATIN SMALL LETTER H WITH HOOK
	`ʘ`: [u8(0x86), 0x42] // U+0298 LATIN LETTER BILABIAL CLICK
	`ǂ`: [u8(0x86), 0x43] // U+01C2 LATIN LETTER ALVEOLAR CLICK
	`ɓ`: [u8(0x86), 0x44] // U+0253 LATIN SMALL LETTER B WITH HOOK
	`ɗ`: [u8(0x86), 0x45] // U+0257 LATIN SMALL LETTER D WITH HOOK
	`ʄ`: [u8(0x86), 0x46] // U+0284 LATIN SMALL LETTER DOTLESS J WITH STROKE AND HOOK
	`ɠ`: [u8(0x86), 0x47] // U+0260 LATIN SMALL LETTER G WITH HOOK
	`Ɠ`: [u8(0x86), 0x48] // U+0193 LATIN CAPITAL LETTER G WITH HOOK
	`œ`: [u8(0x86), 0x49] // U+0153 LATIN SMALL LIGATURE OE
	`Œ`: [u8(0x86), 0x4A] // U+0152 LATIN CAPITAL LIGATURE OE
	`ɨ`: [u8(0x86), 0x4B] // U+0268 LATIN SMALL LETTER I WITH STROKE
	`ʉ`: [u8(0x86), 0x4C] // U+0289 LATIN SMALL LETTER U BAR
	`ɘ`: [u8(0x86), 0x4D] // U+0258 LATIN SMALL LETTER REVERSED E
	`ɵ`: [u8(0x86), 0x4E] // U+0275 LATIN SMALL LETTER BARRED O
	`ə`: [u8(0x86), 0x4F] // U+0259 LATIN SMALL LETTER SCHWA
	`ɜ`: [u8(0x86), 0x50] // U+025C LATIN SMALL LETTER REVERSED OPEN E
	`ɞ`: [u8(0x86), 0x51] // U+025E LATIN SMALL LETTER CLOSED REVERSED OPEN E
	`ɐ`: [u8(0x86), 0x52] // U+0250 LATIN SMALL LETTER TURNED A
	`ɯ`: [u8(0x86), 0x53] // U+026F LATIN SMALL LETTER TURNED M
	`ʊ`: [u8(0x86), 0x54] // U+028A LATIN SMALL LETTER UPSILON
	`ɤ`: [u8(0x86), 0x55] // U+0264 LATIN SMALL LETTER RAMS HORN
	`ʌ`: [u8(0x86), 0x56] // U+028C LATIN SMALL LETTER TURNED V
	`ɔ`: [u8(0x86), 0x57] // U+0254 LATIN SMALL LETTER OPEN O
	`ɑ`: [u8(0x86), 0x58] // U+0251 LATIN SMALL LETTER ALPHA
	`ɒ`: [u8(0x86), 0x59] // U+0252 LATIN SMALL LETTER TURNED ALPHA
	`ʍ`: [u8(0x86), 0x5A] // U+028D LATIN SMALL LETTER TURNED W
	`ɥ`: [u8(0x86), 0x5B] // U+0265 LATIN SMALL LETTER TURNED H
	`ʢ`: [u8(0x86), 0x5C] // U+02A2 LATIN LETTER REVERSED GLOTTAL STOP WITH STROKE
	`ʡ`: [u8(0x86), 0x5D] // U+02A1 LATIN LETTER GLOTTAL STOP WITH STROKE
	`ɕ`: [u8(0x86), 0x5E] // U+0255 LATIN SMALL LETTER C WITH CURL
	`ʑ`: [u8(0x86), 0x5F] // U+0291 LATIN SMALL LETTER Z WITH CURL
	`ɺ`: [u8(0x86), 0x60] // U+027A LATIN SMALL LETTER TURNED R WITH LONG LEG
	`ɧ`: [u8(0x86), 0x61] // U+0267 LATIN SMALL LETTER HENG WITH HOOK
	`ɚ`: [u8(0x86), 0x62] // U+025A LATIN SMALL LETTER SCHWA WITH HOOK
	`ǽ`: [u8(0x86), 0x64] // U+01FD LATIN SMALL LETTER AE WITH ACUTE
	`ὰ`: [u8(0x86), 0x65] // U+1F70 GREEK SMALL LETTER ALPHA WITH VARIA
	`ά`: [u8(0x86), 0x66] // U+1F71 GREEK SMALL LETTER ALPHA WITH OXIA
	`ὲ`: [u8(0x86), 0x6F] // U+1F72 GREEK SMALL LETTER EPSILON WITH VARIA
	`έ`: [u8(0x86), 0x70] // U+1F73 GREEK SMALL LETTER EPSILON WITH OXIA
	`͡`: [u8(0x86), 0x71] // U+0361 COMBINING DOUBLE INVERTED BREVE
	`ˈ`: [u8(0x86), 0x72] // U+02C8 MODIFIER LETTER VERTICAL LINE
	`ˌ`: [u8(0x86), 0x73] // U+02CC MODIFIER LETTER LOW VERTICAL LINE
	`ː`: [u8(0x86), 0x74] // U+02D0 MODIFIER LETTER TRIANGULAR COLON
	`ˑ`: [u8(0x86), 0x75] // U+02D1 MODIFIER LETTER HALF TRIANGULAR COLON
	`̆`: [u8(0x86), 0x76] // U+0306 COMBINING BREVE
	`‿`: [u8(0x86), 0x77] // U+203F UNDERTIE
	`̋`: [u8(0x86), 0x78] // U+030B COMBINING DOUBLE ACUTE ACCENT
	`́`: [u8(0x86), 0x79] // U+0301 COMBINING ACUTE ACCENT
	`̄`: [u8(0x86), 0x7A] // U+0304 COMBINING MACRON
	`̀`: [u8(0x86), 0x7B] // U+0300 COMBINING GRAVE ACCENT
	`̏`: [u8(0x86), 0x7C] // U+030F COMBINING DOUBLE GRAVE ACCENT
	`̌`: [u8(0x86), 0x7D] // U+030C COMBINING CARON
	`̂`: [u8(0x86), 0x7E] // U+0302 COMBINING CIRCUMFLEX ACCENT
	`˥`: [u8(0x86), 0x80] // U+02E5 MODIFIER LETTER EXTRA-HIGH TONE BAR
	`˦`: [u8(0x86), 0x81] // U+02E6 MODIFIER LETTER HIGH TONE BAR
	`˧`: [u8(0x86), 0x82] // U+02E7 MODIFIER LETTER MID TONE BAR
	`˨`: [u8(0x86), 0x83] // U+02E8 MODIFIER LETTER LOW TONE BAR
	`˩`: [u8(0x86), 0x84] // U+02E9 MODIFIER LETTER EXTRA-LOW TONE BAR
	`̥`: [u8(0x86), 0x87] // U+0325 COMBINING RING BELOW
	`̬`: [u8(0x86), 0x88] // U+032C COMBINING CARON BELOW
	`̹`: [u8(0x86), 0x89] // U+0339 COMBINING RIGHT HALF RING BELOW
	`̜`: [u8(0x86), 0x8A] // U+031C COMBINING LEFT HALF RING BELOW
	`̟`: [u8(0x86), 0x8B] // U+031F COMBINING PLUS SIGN BELOW
	`̠`: [u8(0x86), 0x8C] // U+0320 COMBINING MINUS SIGN BELOW
	`̈`: [u8(0x86), 0x8D] // U+0308 COMBINING DIAERESIS
	`̽`: [u8(0x86), 0x8E] // U+033D COMBINING X ABOVE
	`̩`: [u8(0x86), 0x8F] // U+0329 COMBINING VERTICAL LINE BELOW
	`̯`: [u8(0x86), 0x90] // U+032F COMBINING INVERTED BREVE BELOW
	`˞`: [u8(0x86), 0x91] // U+02DE MODIFIER LETTER RHOTIC HOOK
	`̤`: [u8(0x86), 0x92] // U+0324 COMBINING DIAERESIS BELOW
	`̰`: [u8(0x86), 0x93] // U+0330 COMBINING TILDE BELOW
	`̼`: [u8(0x86), 0x94] // U+033C COMBINING SEAGULL BELOW
	`̴`: [u8(0x86), 0x95] // U+0334 COMBINING TILDE OVERLAY
	`̝`: [u8(0x86), 0x96] // U+031D COMBINING UP TACK BELOW
	`̞`: [u8(0x86), 0x97] // U+031E COMBINING DOWN TACK BELOW
	`̘`: [u8(0x86), 0x98] // U+0318 COMBINING LEFT TACK BELOW
	`̙`: [u8(0x86), 0x99] // U+0319 COMBINING RIGHT TACK BELOW
	`̪`: [u8(0x86), 0x9A] // U+032A COMBINING BRIDGE BELOW
	`̺`: [u8(0x86), 0x9B] // U+033A COMBINING INVERTED BRIDGE BELOW
	`̻`: [u8(0x86), 0x9C] // U+033B COMBINING SQUARE BELOW
	`̃`: [u8(0x86), 0x9D] // U+0303 COMBINING TILDE
	`̚`: [u8(0x86), 0x9E] // U+031A COMBINING LEFT ANGLE ABOVE
	`❶`: [u8(0x86), 0x9F] // U+2776 DINGBAT NEGATIVE CIRCLED DIGIT ONE
	`❷`: [u8(0x86), 0xA0] // U+2777 DINGBAT NEGATIVE CIRCLED DIGIT TWO
	`❸`: [u8(0x86), 0xA1] // U+2778 DINGBAT NEGATIVE CIRCLED DIGIT THREE
	`❹`: [u8(0x86), 0xA2] // U+2779 DINGBAT NEGATIVE CIRCLED DIGIT FOUR
	`❺`: [u8(0x86), 0xA3] // U+277A DINGBAT NEGATIVE CIRCLED DIGIT FIVE
	`❻`: [u8(0x86), 0xA4] // U+277B DINGBAT NEGATIVE CIRCLED DIGIT SIX
	`❼`: [u8(0x86), 0xA5] // U+277C DINGBAT NEGATIVE CIRCLED DIGIT SEVEN
	`❽`: [u8(0x86), 0xA6] // U+277D DINGBAT NEGATIVE CIRCLED DIGIT EIGHT
	`❾`: [u8(0x86), 0xA7] // U+277E DINGBAT NEGATIVE CIRCLED DIGIT NINE
	`❿`: [u8(0x86), 0xA8] // U+277F DINGBAT NEGATIVE CIRCLED NUMBER TEN
	`⓫`: [u8(0x86), 0xA9] // U+24EB NEGATIVE CIRCLED NUMBER ELEVEN
	`⓬`: [u8(0x86), 0xAA] // U+24EC NEGATIVE CIRCLED NUMBER TWELVE
	`⓭`: [u8(0x86), 0xAB] // U+24ED NEGATIVE CIRCLED NUMBER THIRTEEN
	`⓮`: [u8(0x86), 0xAC] // U+24EE NEGATIVE CIRCLED NUMBER FOURTEEN
	`⓯`: [u8(0x86), 0xAD] // U+24EF NEGATIVE CIRCLED NUMBER FIFTEEN
	`⓰`: [u8(0x86), 0xAE] // U+24F0 NEGATIVE CIRCLED NUMBER SIXTEEN
	`⓱`: [u8(0x86), 0xAF] // U+24F1 NEGATIVE CIRCLED NUMBER SEVENTEEN
	`⓲`: [u8(0x86), 0xB0] // U+24F2 NEGATIVE CIRCLED NUMBER EIGHTEEN
	`⓳`: [u8(0x86), 0xB1] // U+24F3 NEGATIVE CIRCLED NUMBER NINETEEN
	`⓴`: [u8(0x86), 0xB2] // U+24F4 NEGATIVE CIRCLED NUMBER TWENTY
	`ⅰ`: [u8(0x86), 0xB3] // U+2170 SMALL ROMAN NUMERAL ONE
	`ⅱ`: [u8(0x86), 0xB4] // U+2171 SMALL ROMAN NUMERAL TWO
	`ⅲ`: [u8(0x86), 0xB5] // U+2172 SMALL ROMAN NUMERAL THREE
	`ⅳ`: [u8(0x86), 0xB6] // U+2173 SMALL ROMAN NUMERAL FOUR
	`ⅴ`: [u8(0x86), 0xB7] // U+2174 SMALL ROMAN NUMERAL FIVE
	`ⅵ`: [u8(0x86), 0xB8] // U+2175 SMALL ROMAN NUMERAL SIX
	`ⅶ`: [u8(0x86), 0xB9] // U+2176 SMALL ROMAN NUMERAL SEVEN
	`ⅷ`: [u8(0x86), 0xBA] // U+2177 SMALL ROMAN NUMERAL EIGHT
	`ⅸ`: [u8(0x86), 0xBB] // U+2178 SMALL ROMAN NUMERAL NINE
	`ⅹ`: [u8(0x86), 0xBC] // U+2179 SMALL ROMAN NUMERAL TEN
	`ⅺ`: [u8(0x86), 0xBD] // U+217A SMALL ROMAN NUMERAL ELEVEN
	`ⅻ`: [u8(0x86), 0xBE] // U+217B SMALL ROMAN NUMERAL TWELVE
	`ⓐ`: [u8(0x86), 0xBF] // U+24D0 CIRCLED LATIN SMALL LETTER A
	`ⓑ`: [u8(0x86), 0xC0] // U+24D1 CIRCLED LATIN SMALL LETTER B
	`ⓒ`: [u8(0x86), 0xC1] // U+24D2 CIRCLED LATIN SMALL LETTER C
	`ⓓ`: [u8(0x86), 0xC2] // U+24D3 CIRCLED LATIN SMALL LETTER D
	`ⓔ`: [u8(0x86), 0xC3] // U+24D4 CIRCLED LATIN SMALL LETTER E
	`ⓕ`: [u8(0x86), 0xC4] // U+24D5 CIRCLED LATIN SMALL LETTER F
	`ⓖ`: [u8(0x86), 0xC5] // U+24D6 CIRCLED LATIN SMALL LETTER G
	`ⓗ`: [u8(0x86), 0xC6] // U+24D7 CIRCLED LATIN SMALL LETTER H
	`ⓘ`: [u8(0x86), 0xC7] // U+24D8 CIRCLED LATIN SMALL LETTER I
	`ⓙ`: [u8(0x86), 0xC8] // U+24D9 CIRCLED LATIN SMALL LETTER J
	`ⓚ`: [u8(0x86), 0xC9] // U+24DA CIRCLED LATIN SMALL LETTER K
	`ⓛ`: [u8(0x86), 0xCA] // U+24DB CIRCLED LATIN SMALL LETTER L
	`ⓜ`: [u8(0x86), 0xCB] // U+24DC CIRCLED LATIN SMALL LETTER M
	`ⓝ`: [u8(0x86), 0xCC] // U+24DD CIRCLED LATIN SMALL LETTER N
	`ⓞ`: [u8(0x86), 0xCD] // U+24DE CIRCLED LATIN SMALL LETTER O
	`ⓟ`: [u8(0x86), 0xCE] // U+24DF CIRCLED LATIN SMALL LETTER P
	`ⓠ`: [u8(0x86), 0xCF] // U+24E0 CIRCLED LATIN SMALL LETTER Q
	`ⓡ`: [u8(0x86), 0xD0] // U+24E1 CIRCLED LATIN SMALL LETTER R
	`ⓢ`: [u8(0x86), 0xD1] // U+24E2 CIRCLED LATIN SMALL LETTER S
	`ⓣ`: [u8(0x86), 0xD2] // U+24E3 CIRCLED LATIN SMALL LETTER T
	`ⓤ`: [u8(0x86), 0xD3] // U+24E4 CIRCLED LATIN SMALL LETTER U
	`ⓥ`: [u8(0x86), 0xD4] // U+24E5 CIRCLED LATIN SMALL LETTER V
	`ⓦ`: [u8(0x86), 0xD5] // U+24E6 CIRCLED LATIN SMALL LETTER W
	`ⓧ`: [u8(0x86), 0xD6] // U+24E7 CIRCLED LATIN SMALL LETTER X
	`ⓨ`: [u8(0x86), 0xD7] // U+24E8 CIRCLED LATIN SMALL LETTER Y
	`ⓩ`: [u8(0x86), 0xD8] // U+24E9 CIRCLED LATIN SMALL LETTER Z
	`㋐`: [u8(0x86), 0xD9] // U+32D0 CIRCLED KATAKANA A
	`㋑`: [u8(0x86), 0xDA] // U+32D1 CIRCLED KATAKANA I
	`㋒`: [u8(0x86), 0xDB] // U+32D2 CIRCLED KATAKANA U
	`㋓`: [u8(0x86), 0xDC] // U+32D3 CIRCLED KATAKANA E
	`㋔`: [u8(0x86), 0xDD] // U+32D4 CIRCLED KATAKANA O
	`㋕`: [u8(0x86), 0xDE] // U+32D5 CIRCLED KATAKANA KA
	`㋖`: [u8(0x86), 0xDF] // U+32D6 CIRCLED KATAKANA KI
	`㋗`: [u8(0x86), 0xE0] // U+32D7 CIRCLED KATAKANA KU
	`㋘`: [u8(0x86), 0xE1] // U+32D8 CIRCLED KATAKANA KE
	`㋙`: [u8(0x86), 0xE2] // U+32D9 CIRCLED KATAKANA KO
	`㋚`: [u8(0x86), 0xE3] // U+32DA CIRCLED KATAKANA SA
	`㋛`: [u8(0x86), 0xE4] // U+32DB CIRCLED KATAKANA SI
	`㋜`: [u8(0x86), 0xE5] // U+32DC CIRCLED KATAKANA SU
	`㋝`: [u8(0x86), 0xE6] // U+32DD CIRCLED KATAKANA SE
	`㋞`: [u8(0x86), 0xE7] // U+32DE CIRCLED KATAKANA SO
	`㋟`: [u8(0x86), 0xE8] // U+32DF CIRCLED KATAKANA TA
	`㋠`: [u8(0x86), 0xE9] // U+32E0 CIRCLED KATAKANA TI
	`㋡`: [u8(0x86), 0xEA] // U+32E1 CIRCLED KATAKANA TU
	`㋢`: [u8(0x86), 0xEB] // U+32E2 CIRCLED KATAKANA TE
	`㋣`: [u8(0x86), 0xEC] // U+32E3 CIRCLED KATAKANA TO
	`㋺`: [u8(0x86), 0xED] // U+32FA CIRCLED KATAKANA RO
	`㋩`: [u8(0x86), 0xEE] // U+32E9 CIRCLED KATAKANA HA
	`㋥`: [u8(0x86), 0xEF] // U+32E5 CIRCLED KATAKANA NI
	`㋭`: [u8(0x86), 0xF0] // U+32ED CIRCLED KATAKANA HO
	`㋬`: [u8(0x86), 0xF1] // U+32EC CIRCLED KATAKANA HE
	`⁑`: [u8(0x86), 0xFB] // U+2051 TWO ASTERISKS ALIGNED VERTICALLY
	`⁂`: [u8(0x86), 0xFC] // U+2042 ASTERISM
	`①`: [u8(0x87), 0x40] // U+2460 CIRCLED DIGIT ONE
	`②`: [u8(0x87), 0x41] // U+2461 CIRCLED DIGIT TWO
	`③`: [u8(0x87), 0x42] // U+2462 CIRCLED DIGIT THREE
	`④`: [u8(0x87), 0x43] // U+2463 CIRCLED DIGIT FOUR
	`⑤`: [u8(0x87), 0x44] // U+2464 CIRCLED DIGIT FIVE
	`⑥`: [u8(0x87), 0x45] // U+2465 CIRCLED DIGIT SIX
	`⑦`: [u8(0x87), 0x46] // U+2466 CIRCLED DIGIT SEVEN
	`⑧`: [u8(0x87), 0x47] // U+2467 CIRCLED DIGIT EIGHT
	`⑨`: [u8(0x87), 0x48] // U+2468 CIRCLED DIGIT NINE
	`⑩`: [u8(0x87), 0x49] // U+2469 CIRCLED NUMBER TEN
	`⑪`: [u8(0x87), 0x4A] // U+246A CIRCLED NUMBER ELEVEN
	`⑫`: [u8(0x87), 0x4B] // U+246B CIRCLED NUMBER TWELVE
	`⑬`: [u8(0x87), 0x4C] // U+246C CIRCLED NUMBER THIRTEEN
	`⑭`: [u8(0x87), 0x4D] // U+246D CIRCLED NUMBER FOURTEEN
	`⑮`: [u8(0x87), 0x4E] // U+246E CIRCLED NUMBER FIFTEEN
	`⑯`: [u8(0x87), 0x4F] // U+246F CIRCLED NUMBER SIXTEEN
	`⑰`: [u8(0x87), 0x50] // U+2470 CIRCLED NUMBER SEVENTEEN
	`⑱`: [u8(0x87), 0x51] // U+2471 CIRCLED NUMBER EIGHTEEN
	`⑲`: [u8(0x87), 0x52] // U+2472 CIRCLED NUMBER NINETEEN
	`⑳`: [u8(0x87), 0x53] // U+2473 CIRCLED NUMBER TWENTY
	`Ⅰ`: [u8(0x87), 0x54] // U+2160 ROMAN NUMERAL ONE
	`Ⅱ`: [u8(0x87), 0x55] // U+2161 ROMAN NUMERAL TWO
	`Ⅲ`: [u8(0x87), 0x56] // U+2162 ROMAN NUMERAL THREE
	`Ⅳ`: [u8(0x87), 0x57] // U+2163 ROMAN NUMERAL FOUR
	`Ⅴ`: [u8(0x87), 0x58] // U+2164 ROMAN NUMERAL FIVE
	`Ⅵ`: [u8(0x87), 0x59] // U+2165 ROMAN NUMERAL SIX
	`Ⅶ`: [u8(0x87), 0x5A] // U+2166 ROMAN NUMERAL SEVEN
	`Ⅷ`: [u8(0x87), 0x5B] // U+2167 ROMAN NUMERAL EIGHT
	`Ⅸ`: [u8(0x87), 0x5C] // U+2168 ROMAN NUMERAL NINE
	`Ⅹ`: [u8(0x87), 0x5D] // U+2169 ROMAN NUMERAL TEN
	`Ⅺ`: [u8(0x87), 0x5E] // U+216A ROMAN NUMERAL ELEVEN
	`㍉`: [u8(0x87), 0x5F] // U+3349 SQUARE MIRI
	`㌔`: [u8(0x87), 0x60] // U+3314 SQUARE KIRO
	`㌢`: [u8(0x87), 0x61] // U+3322 SQUARE SENTI
	`㍍`: [u8(0x87), 0x62] // U+334D SQUARE MEETORU
	`㌘`: [u8(0x87), 0x63] // U+3318 SQUARE GURAMU
	`㌧`: [u8(0x87), 0x64] // U+3327 SQUARE TON
	`㌃`: [u8(0x87), 0x65] // U+3303 SQUARE AARU
	`㌶`: [u8(0x87), 0x66] // U+3336 SQUARE HEKUTAARU
	`㍑`: [u8(0x87), 0x67] // U+3351 SQUARE RITTORU
	`㍗`: [u8(0x87), 0x68] // U+3357 SQUARE WATTO
	`㌍`: [u8(0x87), 0x69] // U+330D SQUARE KARORII
	`㌦`: [u8(0x87), 0x6A] // U+3326 SQUARE DORU
	`㌣`: [u8(0x87), 0x6B] // U+3323 SQUARE SENTO
	`㌫`: [u8(0x87), 0x6C] // U+332B SQUARE PAASENTO
	`㍊`: [u8(0x87), 0x6D] // U+334A SQUARE MIRIBAARU
	`㌻`: [u8(0x87), 0x6E] // U+333B SQUARE PEEZI
	`㎜`: [u8(0x87), 0x6F] // U+339C SQUARE MM
	`㎝`: [u8(0x87), 0x70] // U+339D SQUARE CM
	`㎞`: [u8(0x87), 0x71] // U+339E SQUARE KM
	`㎎`: [u8(0x87), 0x72] // U+338E SQUARE MG
	`㎏`: [u8(0x87), 0x73] // U+338F SQUARE KG
	`㏄`: [u8(0x87), 0x74] // U+33C4 SQUARE CC
	`㎡`: [u8(0x87), 0x75] // U+33A1 SQUARE M SQUARED
	`Ⅻ`: [u8(0x87), 0x76] // U+216B ROMAN NUMERAL TWELVE
	`㍻`: [u8(0x87), 0x7E] // U+337B SQUARE ERA NAME HEISEI
	`〝`: [u8(0x87), 0x80] // U+301D REVERSED DOUBLE PRIME QUOTATION MARK
	`〟`: [u8(0x87), 0x81] // U+301F LOW DOUBLE PRIME QUOTATION MARK
	`№`: [u8(0x87), 0x82] // U+2116 NUMERO SIGN
	`㏍`: [u8(0x87), 0x83] // U+33CD SQUARE KK
	`℡`: [u8(0x87), 0x84] // U+2121 TELEPHONE SIGN
	`㊤`: [u8(0x87), 0x85] // U+32A4 CIRCLED IDEOGRAPH HIGH
	`㊥`: [u8(0x87), 0x86] // U+32A5 CIRCLED IDEOGRAPH CENTRE
	`㊦`: [u8(0x87), 0x87] // U+32A6 CIRCLED IDEOGRAPH LOW
	`㊧`: [u8(0x87), 0x88] // U+32A7 CIRCLED IDEOGRAPH LEFT
	`㊨`: [u8(0x87), 0x89] // U+32A8 CIRCLED IDEOGRAPH RIGHT
	`㈱`: [u8(0x87), 0x8A] // U+3231 PARENTHESIZED IDEOGRAPH STOCK
	`㈲`: [u8(0x87), 0x8B] // U+3232 PARENTHESIZED IDEOGRAPH HAVE
	`㈹`: [u8(0x87), 0x8C] // U+3239 PARENTHESIZED IDEOGRAPH REPRESENT
	`㍾`: [u8(0x87), 0x8D] // U+337E SQUARE ERA NAME MEIZI
	`㍽`: [u8(0x87), 0x8E] // U+337D SQUARE ERA NAME TAISYOU
	`㍼`: [u8(0x87), 0x8F] // U+337C SQUARE ERA NAME SYOUWA
	`∮`: [u8(0x87), 0x93] // U+222E CONTOUR INTEGRAL
	`∟`: [u8(0x87), 0x98] // U+221F RIGHT ANGLE
	`⊿`: [u8(0x87), 0x99] // U+22BF RIGHT TRIANGLE
	`❖`: [u8(0x87), 0x9D] // U+2756 BLACK DIAMOND MINUS WHITE X
	`☞`: [u8(0x87), 0x9E] // U+261E WHITE RIGHT POINTING INDEX
	`俱`: [u8(0x87), 0x9F] // U+4FF1 <cjk>
	`𠀋`: [u8(0x87), 0xA0] // U+2000B <cjk>
	`㐂`: [u8(0x87), 0xA1] // U+3402 <cjk>
	`丨`: [u8(0x87), 0xA2] // U+4E28 <cjk>
	`丯`: [u8(0x87), 0xA3] // U+4E2F <cjk>
	`丰`: [u8(0x87), 0xA4] // U+4E30 <cjk>
	`亍`: [u8(0x87), 0xA5] // U+4E8D <cjk>
	`仡`: [u8(0x87), 0xA6] // U+4EE1 <cjk>
	`份`: [u8(0x87), 0xA7] // U+4EFD <cjk>
	`仿`: [u8(0x87), 0xA8] // U+4EFF <cjk>
	`伃`: [u8(0x87), 0xA9] // U+4F03 <cjk>
	`伋`: [u8(0x87), 0xAA] // U+4F0B <cjk>
	`你`: [u8(0x87), 0xAB] // U+4F60 <cjk>
	`佈`: [u8(0x87), 0xAC] // U+4F48 <cjk>
	`佉`: [u8(0x87), 0xAD] // U+4F49 <cjk>
	`佖`: [u8(0x87), 0xAE] // U+4F56 <cjk>
	`佟`: [u8(0x87), 0xAF] // U+4F5F <cjk>
	`佪`: [u8(0x87), 0xB0] // U+4F6A <cjk>
	`佬`: [u8(0x87), 0xB1] // U+4F6C <cjk>
	`佾`: [u8(0x87), 0xB2] // U+4F7E <cjk>
	`侊`: [u8(0x87), 0xB3] // U+4F8A <cjk>
	`侔`: [u8(0x87), 0xB4] // U+4F94 <cjk>
	`侗`: [u8(0x87), 0xB5] // U+4F97 <cjk>
	`侮`: [u8(0x87), 0xB6] // U+FA30 CJK COMPATIBILITY IDEOGRAPH-FA30
	`俉`: [u8(0x87), 0xB7] // U+4FC9 <cjk>
	`俠`: [u8(0x87), 0xB8] // U+4FE0 <cjk>
	`倁`: [u8(0x87), 0xB9] // U+5001 <cjk>
	`倂`: [u8(0x87), 0xBA] // U+5002 <cjk>
	`倎`: [u8(0x87), 0xBB] // U+500E <cjk>
	`倘`: [u8(0x87), 0xBC] // U+5018 <cjk>
	`倧`: [u8(0x87), 0xBD] // U+5027 <cjk>
	`倮`: [u8(0x87), 0xBE] // U+502E <cjk>
	`偀`: [u8(0x87), 0xBF] // U+5040 <cjk>
	`倻`: [u8(0x87), 0xC0] // U+503B <cjk>
	`偁`: [u8(0x87), 0xC1] // U+5041 <cjk>
	`傔`: [u8(0x87), 0xC2] // U+5094 <cjk>
	`僌`: [u8(0x87), 0xC3] // U+50CC <cjk>
	`僲`: [u8(0x87), 0xC4] // U+50F2 <cjk>
	`僐`: [u8(0x87), 0xC5] // U+50D0 <cjk>
	`僦`: [u8(0x87), 0xC6] // U+50E6 <cjk>
	`僧`: [u8(0x87), 0xC7] // U+FA31 CJK COMPATIBILITY IDEOGRAPH-FA31
	`儆`: [u8(0x87), 0xC8] // U+5106 <cjk>
	`儃`: [u8(0x87), 0xC9] // U+5103 <cjk>
	`儋`: [u8(0x87), 0xCA] // U+510B <cjk>
	`儞`: [u8(0x87), 0xCB] // U+511E <cjk>
	`儵`: [u8(0x87), 0xCC] // U+5135 <cjk>
	`兊`: [u8(0x87), 0xCD] // U+514A <cjk>
	`免`: [u8(0x87), 0xCE] // U+FA32 CJK COMPATIBILITY IDEOGRAPH-FA32
	`兕`: [u8(0x87), 0xCF] // U+5155 <cjk>
	`兗`: [u8(0x87), 0xD0] // U+5157 <cjk>
	`㒵`: [u8(0x87), 0xD1] // U+34B5 <cjk>
	`冝`: [u8(0x87), 0xD2] // U+519D <cjk>
	`凃`: [u8(0x87), 0xD3] // U+51C3 <cjk>
	`凊`: [u8(0x87), 0xD4] // U+51CA <cjk>
	`凞`: [u8(0x87), 0xD5] // U+51DE <cjk>
	`凢`: [u8(0x87), 0xD6] // U+51E2 <cjk>
	`凮`: [u8(0x87), 0xD7] // U+51EE <cjk>
	`刁`: [u8(0x87), 0xD8] // U+5201 <cjk>
	`㓛`: [u8(0x87), 0xD9] // U+34DB <cjk>
	`刓`: [u8(0x87), 0xDA] // U+5213 <cjk>
	`刕`: [u8(0x87), 0xDB] // U+5215 <cjk>
	`剉`: [u8(0x87), 0xDC] // U+5249 <cjk>
	`剗`: [u8(0x87), 0xDD] // U+5257 <cjk>
	`剡`: [u8(0x87), 0xDE] // U+5261 <cjk>
	`劓`: [u8(0x87), 0xDF] // U+5293 <cjk>
	`勈`: [u8(0x87), 0xE0] // U+52C8 <cjk>
	`勉`: [u8(0x87), 0xE1] // U+FA33 CJK COMPATIBILITY IDEOGRAPH-FA33
	`勌`: [u8(0x87), 0xE2] // U+52CC <cjk>
	`勐`: [u8(0x87), 0xE3] // U+52D0 <cjk>
	`勖`: [u8(0x87), 0xE4] // U+52D6 <cjk>
	`勛`: [u8(0x87), 0xE5] // U+52DB <cjk>
	`勤`: [u8(0x87), 0xE6] // U+FA34 CJK COMPATIBILITY IDEOGRAPH-FA34
	`勰`: [u8(0x87), 0xE7] // U+52F0 <cjk>
	`勻`: [u8(0x87), 0xE8] // U+52FB <cjk>
	`匀`: [u8(0x87), 0xE9] // U+5300 <cjk>
	`匇`: [u8(0x87), 0xEA] // U+5307 <cjk>
	`匜`: [u8(0x87), 0xEB] // U+531C <cjk>
	`卑`: [u8(0x87), 0xEC] // U+FA35 CJK COMPATIBILITY IDEOGRAPH-FA35
	`卡`: [u8(0x87), 0xED] // U+5361 <cjk>
	`卣`: [u8(0x87), 0xEE] // U+5363 <cjk>
	`卽`: [u8(0x87), 0xEF] // U+537D <cjk>
	`厓`: [u8(0x87), 0xF0] // U+5393 <cjk>
	`厝`: [u8(0x87), 0xF1] // U+539D <cjk>
	`厲`: [u8(0x87), 0xF2] // U+53B2 <cjk>
	`吒`: [u8(0x87), 0xF3] // U+5412 <cjk>
	`吧`: [u8(0x87), 0xF4] // U+5427 <cjk>
	`呍`: [u8(0x87), 0xF5] // U+544D <cjk>
	`咜`: [u8(0x87), 0xF6] // U+549C <cjk>
	`呫`: [u8(0x87), 0xF7] // U+546B <cjk>
	`呴`: [u8(0x87), 0xF8] // U+5474 <cjk>
	`呿`: [u8(0x87), 0xF9] // U+547F <cjk>
	`咈`: [u8(0x87), 0xFA] // U+5488 <cjk>
	`咖`: [u8(0x87), 0xFB] // U+5496 <cjk>
	`咡`: [u8(0x87), 0xFC] // U+54A1 <cjk>
	`咩`: [u8(0x88), 0x40] // U+54A9 <cjk>
	`哆`: [u8(0x88), 0x41] // U+54C6 <cjk>
	`哿`: [u8(0x88), 0x42] // U+54FF <cjk>
	`唎`: [u8(0x88), 0x43] // U+550E <cjk>
	`唫`: [u8(0x88), 0x44] // U+552B <cjk>
	`唵`: [u8(0x88), 0x45] // U+5535 <cjk>
	`啐`: [u8(0x88), 0x46] // U+5550 <cjk>
	`啞`: [u8(0x88), 0x47] // U+555E <cjk>
	`喁`: [u8(0x88), 0x48] // U+5581 <cjk>
	`喆`: [u8(0x88), 0x49] // U+5586 <cjk>
	`喎`: [u8(0x88), 0x4A] // U+558E <cjk>
	`喝`: [u8(0x88), 0x4B] // U+FA36 CJK COMPATIBILITY IDEOGRAPH-FA36
	`喭`: [u8(0x88), 0x4C] // U+55AD <cjk>
	`嗎`: [u8(0x88), 0x4D] // U+55CE <cjk>
	`嘆`: [u8(0x88), 0x4E] // U+FA37 CJK COMPATIBILITY IDEOGRAPH-FA37
	`嘈`: [u8(0x88), 0x4F] // U+5608 <cjk>
	`嘎`: [u8(0x88), 0x50] // U+560E <cjk>
	`嘻`: [u8(0x88), 0x51] // U+563B <cjk>
	`噉`: [u8(0x88), 0x52] // U+5649 <cjk>
	`噶`: [u8(0x88), 0x53] // U+5676 <cjk>
	`噦`: [u8(0x88), 0x54] // U+5666 <cjk>
	`器`: [u8(0x88), 0x55] // U+FA38 CJK COMPATIBILITY IDEOGRAPH-FA38
	`噯`: [u8(0x88), 0x56] // U+566F <cjk>
	`噱`: [u8(0x88), 0x57] // U+5671 <cjk>
	`噲`: [u8(0x88), 0x58] // U+5672 <cjk>
	`嚙`: [u8(0x88), 0x59] // U+5699 <cjk>
	`嚞`: [u8(0x88), 0x5A] // U+569E <cjk>
	`嚩`: [u8(0x88), 0x5B] // U+56A9 <cjk>
	`嚬`: [u8(0x88), 0x5C] // U+56AC <cjk>
	`嚳`: [u8(0x88), 0x5D] // U+56B3 <cjk>
	`囉`: [u8(0x88), 0x5E] // U+56C9 <cjk>
	`囊`: [u8(0x88), 0x5F] // U+56CA <cjk>
	`圊`: [u8(0x88), 0x60] // U+570A <cjk>
	`𡈽`: [u8(0x88), 0x61] // U+2123D <cjk>
	`圡`: [u8(0x88), 0x62] // U+5721 <cjk>
	`圯`: [u8(0x88), 0x63] // U+572F <cjk>
	`圳`: [u8(0x88), 0x64] // U+5733 <cjk>
	`圴`: [u8(0x88), 0x65] // U+5734 <cjk>
	`坰`: [u8(0x88), 0x66] // U+5770 <cjk>
	`坷`: [u8(0x88), 0x67] // U+5777 <cjk>
	`坼`: [u8(0x88), 0x68] // U+577C <cjk>
	`垜`: [u8(0x88), 0x69] // U+579C <cjk>
	`﨏`: [u8(0x88), 0x6A] // U+FA0F CJK COMPATIBILITY IDEOGRAPH-FA0F
	`𡌛`: [u8(0x88), 0x6B] // U+2131B <cjk>
	`垸`: [u8(0x88), 0x6C] // U+57B8 <cjk>
	`埇`: [u8(0x88), 0x6D] // U+57C7 <cjk>
	`埈`: [u8(0x88), 0x6E] // U+57C8 <cjk>
	`埏`: [u8(0x88), 0x6F] // U+57CF <cjk>
	`埤`: [u8(0x88), 0x70] // U+57E4 <cjk>
	`埭`: [u8(0x88), 0x71] // U+57ED <cjk>
	`埵`: [u8(0x88), 0x72] // U+57F5 <cjk>
	`埶`: [u8(0x88), 0x73] // U+57F6 <cjk>
	`埿`: [u8(0x88), 0x74] // U+57FF <cjk>
	`堉`: [u8(0x88), 0x75] // U+5809 <cjk>
	`塚`: [u8(0x88), 0x76] // U+FA10 CJK COMPATIBILITY IDEOGRAPH-FA10
	`塡`: [u8(0x88), 0x77] // U+5861 <cjk>
	`塤`: [u8(0x88), 0x78] // U+5864 <cjk>
	`塀`: [u8(0x88), 0x79] // U+FA39 CJK COMPATIBILITY IDEOGRAPH-FA39
	`塼`: [u8(0x88), 0x7A] // U+587C <cjk>
	`墉`: [u8(0x88), 0x7B] // U+5889 <cjk>
	`增`: [u8(0x88), 0x7C] // U+589E <cjk>
	`墨`: [u8(0x88), 0x7D] // U+FA3A CJK COMPATIBILITY IDEOGRAPH-FA3A
	`墩`: [u8(0x88), 0x7E] // U+58A9 <cjk>
	`𡑮`: [u8(0x88), 0x80] // U+2146E <cjk>
	`壒`: [u8(0x88), 0x81] // U+58D2 <cjk>
	`壎`: [u8(0x88), 0x82] // U+58CE <cjk>
	`壔`: [u8(0x88), 0x83] // U+58D4 <cjk>
	`壚`: [u8(0x88), 0x84] // U+58DA <cjk>
	`壠`: [u8(0x88), 0x85] // U+58E0 <cjk>
	`壩`: [u8(0x88), 0x86] // U+58E9 <cjk>
	`夌`: [u8(0x88), 0x87] // U+590C <cjk>
	`虁`: [u8(0x88), 0x88] // U+8641 <cjk>
	`奝`: [u8(0x88), 0x89] // U+595D <cjk>
	`奭`: [u8(0x88), 0x8A] // U+596D <cjk>
	`妋`: [u8(0x88), 0x8B] // U+598B <cjk>
	`妒`: [u8(0x88), 0x8C] // U+5992 <cjk>
	`妤`: [u8(0x88), 0x8D] // U+59A4 <cjk>
	`姃`: [u8(0x88), 0x8E] // U+59C3 <cjk>
	`姒`: [u8(0x88), 0x8F] // U+59D2 <cjk>
	`姝`: [u8(0x88), 0x90] // U+59DD <cjk>
	`娓`: [u8(0x88), 0x91] // U+5A13 <cjk>
	`娣`: [u8(0x88), 0x92] // U+5A23 <cjk>
	`婧`: [u8(0x88), 0x93] // U+5A67 <cjk>
	`婭`: [u8(0x88), 0x94] // U+5A6D <cjk>
	`婷`: [u8(0x88), 0x95] // U+5A77 <cjk>
	`婾`: [u8(0x88), 0x96] // U+5A7E <cjk>
	`媄`: [u8(0x88), 0x97] // U+5A84 <cjk>
	`媞`: [u8(0x88), 0x98] // U+5A9E <cjk>
	`媧`: [u8(0x88), 0x99] // U+5AA7 <cjk>
	`嫄`: [u8(0x88), 0x9A] // U+5AC4 <cjk>
	`𡢽`: [u8(0x88), 0x9B] // U+218BD <cjk>
	`嬙`: [u8(0x88), 0x9C] // U+5B19 <cjk>
	`嬥`: [u8(0x88), 0x9D] // U+5B25 <cjk>
	`剝`: [u8(0x88), 0x9E] // U+525D <cjk>
	`亜`: [u8(0x88), 0x9F] // U+4E9C <cjk>
	`唖`: [u8(0x88), 0xA0] // U+5516 <cjk>
	`娃`: [u8(0x88), 0xA1] // U+5A03 <cjk>
	`阿`: [u8(0x88), 0xA2] // U+963F <cjk>
	`哀`: [u8(0x88), 0xA3] // U+54C0 <cjk>
	`愛`: [u8(0x88), 0xA4] // U+611B <cjk>
	`挨`: [u8(0x88), 0xA5] // U+6328 <cjk>
	`姶`: [u8(0x88), 0xA6] // U+59F6 <cjk>
	`逢`: [u8(0x88), 0xA7] // U+9022 <cjk>
	`葵`: [u8(0x88), 0xA8] // U+8475 <cjk>
	`茜`: [u8(0x88), 0xA9] // U+831C <cjk>
	`穐`: [u8(0x88), 0xAA] // U+7A50 <cjk>
	`悪`: [u8(0x88), 0xAB] // U+60AA <cjk>
	`握`: [u8(0x88), 0xAC] // U+63E1 <cjk>
	`渥`: [u8(0x88), 0xAD] // U+6E25 <cjk>
	`旭`: [u8(0x88), 0xAE] // U+65ED <cjk>
	`葦`: [u8(0x88), 0xAF] // U+8466 <cjk>
	`芦`: [u8(0x88), 0xB0] // U+82A6 <cjk>
	`鯵`: [u8(0x88), 0xB1] // U+9BF5 <cjk>
	`梓`: [u8(0x88), 0xB2] // U+6893 <cjk>
	`圧`: [u8(0x88), 0xB3] // U+5727 <cjk>
	`斡`: [u8(0x88), 0xB4] // U+65A1 <cjk>
	`扱`: [u8(0x88), 0xB5] // U+6271 <cjk>
	`宛`: [u8(0x88), 0xB6] // U+5B9B <cjk>
	`姐`: [u8(0x88), 0xB7] // U+59D0 <cjk>
	`虻`: [u8(0x88), 0xB8] // U+867B <cjk>
	`飴`: [u8(0x88), 0xB9] // U+98F4 <cjk>
	`絢`: [u8(0x88), 0xBA] // U+7D62 <cjk>
	`綾`: [u8(0x88), 0xBB] // U+7DBE <cjk>
	`鮎`: [u8(0x88), 0xBC] // U+9B8E <cjk>
	`或`: [u8(0x88), 0xBD] // U+6216 <cjk>
	`粟`: [u8(0x88), 0xBE] // U+7C9F <cjk>
	`袷`: [u8(0x88), 0xBF] // U+88B7 <cjk>
	`安`: [u8(0x88), 0xC0] // U+5B89 <cjk>
	`庵`: [u8(0x88), 0xC1] // U+5EB5 <cjk>
	`按`: [u8(0x88), 0xC2] // U+6309 <cjk>
	`暗`: [u8(0x88), 0xC3] // U+6697 <cjk>
	`案`: [u8(0x88), 0xC4] // U+6848 <cjk>
	`闇`: [u8(0x88), 0xC5] // U+95C7 <cjk>
	`鞍`: [u8(0x88), 0xC6] // U+978D <cjk>
	`杏`: [u8(0x88), 0xC7] // U+674F <cjk>
	`以`: [u8(0x88), 0xC8] // U+4EE5 <cjk>
	`伊`: [u8(0x88), 0xC9] // U+4F0A <cjk>
	`位`: [u8(0x88), 0xCA] // U+4F4D <cjk>
	`依`: [u8(0x88), 0xCB] // U+4F9D <cjk>
	`偉`: [u8(0x88), 0xCC] // U+5049 <cjk>
	`囲`: [u8(0x88), 0xCD] // U+56F2 <cjk>
	`夷`: [u8(0x88), 0xCE] // U+5937 <cjk>
	`委`: [u8(0x88), 0xCF] // U+59D4 <cjk>
	`威`: [u8(0x88), 0xD0] // U+5A01 <cjk>
	`尉`: [u8(0x88), 0xD1] // U+5C09 <cjk>
	`惟`: [u8(0x88), 0xD2] // U+60DF <cjk>
	`意`: [u8(0x88), 0xD3] // U+610F <cjk>
	`慰`: [u8(0x88), 0xD4] // U+6170 <cjk>
	`易`: [u8(0x88), 0xD5] // U+6613 <cjk>
	`椅`: [u8(0x88), 0xD6] // U+6905 <cjk>
	`為`: [u8(0x88), 0xD7] // U+70BA <cjk>
	`畏`: [u8(0x88), 0xD8] // U+754F <cjk>
	`異`: [u8(0x88), 0xD9] // U+7570 <cjk>
	`移`: [u8(0x88), 0xDA] // U+79FB <cjk>
	`維`: [u8(0x88), 0xDB] // U+7DAD <cjk>
	`緯`: [u8(0x88), 0xDC] // U+7DEF <cjk>
	`胃`: [u8(0x88), 0xDD] // U+80C3 <cjk>
	`萎`: [u8(0x88), 0xDE] // U+840E <cjk>
	`衣`: [u8(0x88), 0xDF] // U+8863 <cjk>
	`謂`: [u8(0x88), 0xE0] // U+8B02 <cjk>
	`違`: [u8(0x88), 0xE1] // U+9055 <cjk>
	`遺`: [u8(0x88), 0xE2] // U+907A <cjk>
	`医`: [u8(0x88), 0xE3] // U+533B <cjk>
	`井`: [u8(0x88), 0xE4] // U+4E95 <cjk>
	`亥`: [u8(0x88), 0xE5] // U+4EA5 <cjk>
	`域`: [u8(0x88), 0xE6] // U+57DF <cjk>
	`育`: [u8(0x88), 0xE7] // U+80B2 <cjk>
	`郁`: [u8(0x88), 0xE8] // U+90C1 <cjk>
	`磯`: [u8(0x88), 0xE9] // U+78EF <cjk>
	`一`: [u8(0x88), 0xEA] // U+4E00 <cjk>
	`壱`: [u8(0x88), 0xEB] // U+58F1 <cjk>
	`溢`: [u8(0x88), 0xEC] // U+6EA2 <cjk>
	`逸`: [u8(0x88), 0xED] // U+9038 <cjk>
	`稲`: [u8(0x88), 0xEE] // U+7A32 <cjk>
	`茨`: [u8(0x88), 0xEF] // U+8328 <cjk>
	`芋`: [u8(0x88), 0xF0] // U+828B <cjk>
	`鰯`: [u8(0x88), 0xF1] // U+9C2F <cjk>
	`允`: [u8(0x88), 0xF2] // U+5141 <cjk>
	`印`: [u8(0x88), 0xF3] // U+5370 <cjk>
	`咽`: [u8(0x88), 0xF4] // U+54BD <cjk>
	`員`: [u8(0x88), 0xF5] // U+54E1 <cjk>
	`因`: [u8(0x88), 0xF6] // U+56E0 <cjk>
	`姻`: [u8(0x88), 0xF7] // U+59FB <cjk>
	`引`: [u8(0x88), 0xF8] // U+5F15 <cjk>
	`飲`: [u8(0x88), 0xF9] // U+98F2 <cjk>
	`淫`: [u8(0x88), 0xFA] // U+6DEB <cjk>
	`胤`: [u8(0x88), 0xFB] // U+80E4 <cjk>
	`蔭`: [u8(0x88), 0xFC] // U+852D <cjk>
	`院`: [u8(0x89), 0x40] // U+9662 <cjk>
	`陰`: [u8(0x89), 0x41] // U+9670 <cjk>
	`隠`: [u8(0x89), 0x42] // U+96A0 <cjk>
	`韻`: [u8(0x89), 0x43] // U+97FB <cjk>
	`吋`: [u8(0x89), 0x44] // U+540B <cjk>
	`右`: [u8(0x89), 0x45] // U+53F3 <cjk>
	`宇`: [u8(0x89), 0x46] // U+5B87 <cjk>
	`烏`: [u8(0x89), 0x47] // U+70CF <cjk>
	`羽`: [u8(0x89), 0x48] // U+7FBD <cjk>
	`迂`: [u8(0x89), 0x49] // U+8FC2 <cjk>
	`雨`: [u8(0x89), 0x4A] // U+96E8 <cjk>
	`卯`: [u8(0x89), 0x4B] // U+536F <cjk>
	`鵜`: [u8(0x89), 0x4C] // U+9D5C <cjk>
	`窺`: [u8(0x89), 0x4D] // U+7ABA <cjk>
	`丑`: [u8(0x89), 0x4E] // U+4E11 <cjk>
	`碓`: [u8(0x89), 0x4F] // U+7893 <cjk>
	`臼`: [u8(0x89), 0x50] // U+81FC <cjk>
	`渦`: [u8(0x89), 0x51] // U+6E26 <cjk>
	`嘘`: [u8(0x89), 0x52] // U+5618 <cjk>
	`唄`: [u8(0x89), 0x53] // U+5504 <cjk>
	`欝`: [u8(0x89), 0x54] // U+6B1D <cjk>
	`蔚`: [u8(0x89), 0x55] // U+851A <cjk>
	`鰻`: [u8(0x89), 0x56] // U+9C3B <cjk>
	`姥`: [u8(0x89), 0x57] // U+59E5 <cjk>
	`厩`: [u8(0x89), 0x58] // U+53A9 <cjk>
	`浦`: [u8(0x89), 0x59] // U+6D66 <cjk>
	`瓜`: [u8(0x89), 0x5A] // U+74DC <cjk>
	`閏`: [u8(0x89), 0x5B] // U+958F <cjk>
	`噂`: [u8(0x89), 0x5C] // U+5642 <cjk>
	`云`: [u8(0x89), 0x5D] // U+4E91 <cjk>
	`運`: [u8(0x89), 0x5E] // U+904B <cjk>
	`雲`: [u8(0x89), 0x5F] // U+96F2 <cjk>
	`荏`: [u8(0x89), 0x60] // U+834F <cjk>
	`餌`: [u8(0x89), 0x61] // U+990C <cjk>
	`叡`: [u8(0x89), 0x62] // U+53E1 <cjk>
	`営`: [u8(0x89), 0x63] // U+55B6 <cjk>
	`嬰`: [u8(0x89), 0x64] // U+5B30 <cjk>
	`影`: [u8(0x89), 0x65] // U+5F71 <cjk>
	`映`: [u8(0x89), 0x66] // U+6620 <cjk>
	`曳`: [u8(0x89), 0x67] // U+66F3 <cjk>
	`栄`: [u8(0x89), 0x68] // U+6804 <cjk>
	`永`: [u8(0x89), 0x69] // U+6C38 <cjk>
	`泳`: [u8(0x89), 0x6A] // U+6CF3 <cjk>
	`洩`: [u8(0x89), 0x6B] // U+6D29 <cjk>
	`瑛`: [u8(0x89), 0x6C] // U+745B <cjk>
	`盈`: [u8(0x89), 0x6D] // U+76C8 <cjk>
	`穎`: [u8(0x89), 0x6E] // U+7A4E <cjk>
	`頴`: [u8(0x89), 0x6F] // U+9834 <cjk>
	`英`: [u8(0x89), 0x70] // U+82F1 <cjk>
	`衛`: [u8(0x89), 0x71] // U+885B <cjk>
	`詠`: [u8(0x89), 0x72] // U+8A60 <cjk>
	`鋭`: [u8(0x89), 0x73] // U+92ED <cjk>
	`液`: [u8(0x89), 0x74] // U+6DB2 <cjk>
	`疫`: [u8(0x89), 0x75] // U+75AB <cjk>
	`益`: [u8(0x89), 0x76] // U+76CA <cjk>
	`駅`: [u8(0x89), 0x77] // U+99C5 <cjk>
	`悦`: [u8(0x89), 0x78] // U+60A6 <cjk>
	`謁`: [u8(0x89), 0x79] // U+8B01 <cjk>
	`越`: [u8(0x89), 0x7A] // U+8D8A <cjk>
	`閲`: [u8(0x89), 0x7B] // U+95B2 <cjk>
	`榎`: [u8(0x89), 0x7C] // U+698E <cjk>
	`厭`: [u8(0x89), 0x7D] // U+53AD <cjk>
	`円`: [u8(0x89), 0x7E] // U+5186 <cjk>
	`園`: [u8(0x89), 0x80] // U+5712 <cjk>
	`堰`: [u8(0x89), 0x81] // U+5830 <cjk>
	`奄`: [u8(0x89), 0x82] // U+5944 <cjk>
	`宴`: [u8(0x89), 0x83] // U+5BB4 <cjk>
	`延`: [u8(0x89), 0x84] // U+5EF6 <cjk>
	`怨`: [u8(0x89), 0x85] // U+6028 <cjk>
	`掩`: [u8(0x89), 0x86] // U+63A9 <cjk>
	`援`: [u8(0x89), 0x87] // U+63F4 <cjk>
	`沿`: [u8(0x89), 0x88] // U+6CBF <cjk>
	`演`: [u8(0x89), 0x89] // U+6F14 <cjk>
	`炎`: [u8(0x89), 0x8A] // U+708E <cjk>
	`焔`: [u8(0x89), 0x8B] // U+7114 <cjk>
	`煙`: [u8(0x89), 0x8C] // U+7159 <cjk>
	`燕`: [u8(0x89), 0x8D] // U+71D5 <cjk>
	`猿`: [u8(0x89), 0x8E] // U+733F <cjk>
	`縁`: [u8(0x89), 0x8F] // U+7E01 <cjk>
	`艶`: [u8(0x89), 0x90] // U+8276 <cjk>
	`苑`: [u8(0x89), 0x91] // U+82D1 <cjk>
	`薗`: [u8(0x89), 0x92] // U+8597 <cjk>
	`遠`: [u8(0x89), 0x93] // U+9060 <cjk>
	`鉛`: [u8(0x89), 0x94] // U+925B <cjk>
	`鴛`: [u8(0x89), 0x95] // U+9D1B <cjk>
	`塩`: [u8(0x89), 0x96] // U+5869 <cjk>
	`於`: [u8(0x89), 0x97] // U+65BC <cjk>
	`汚`: [u8(0x89), 0x98] // U+6C5A <cjk>
	`甥`: [u8(0x89), 0x99] // U+7525 <cjk>
	`凹`: [u8(0x89), 0x9A] // U+51F9 <cjk>
	`央`: [u8(0x89), 0x9B] // U+592E <cjk>
	`奥`: [u8(0x89), 0x9C] // U+5965 <cjk>
	`往`: [u8(0x89), 0x9D] // U+5F80 <cjk>
	`応`: [u8(0x89), 0x9E] // U+5FDC <cjk>
	`押`: [u8(0x89), 0x9F] // U+62BC <cjk>
	`旺`: [u8(0x89), 0xA0] // U+65FA <cjk>
	`横`: [u8(0x89), 0xA1] // U+6A2A <cjk>
	`欧`: [u8(0x89), 0xA2] // U+6B27 <cjk>
	`殴`: [u8(0x89), 0xA3] // U+6BB4 <cjk>
	`王`: [u8(0x89), 0xA4] // U+738B <cjk>
	`翁`: [u8(0x89), 0xA5] // U+7FC1 <cjk>
	`襖`: [u8(0x89), 0xA6] // U+8956 <cjk>
	`鴬`: [u8(0x89), 0xA7] // U+9D2C <cjk>
	`鴎`: [u8(0x89), 0xA8] // U+9D0E <cjk>
	`黄`: [u8(0x89), 0xA9] // U+9EC4 <cjk>
	`岡`: [u8(0x89), 0xAA] // U+5CA1 <cjk>
	`沖`: [u8(0x89), 0xAB] // U+6C96 <cjk>
	`荻`: [u8(0x89), 0xAC] // U+837B <cjk>
	`億`: [u8(0x89), 0xAD] // U+5104 <cjk>
	`屋`: [u8(0x89), 0xAE] // U+5C4B <cjk>
	`憶`: [u8(0x89), 0xAF] // U+61B6 <cjk>
	`臆`: [u8(0x89), 0xB0] // U+81C6 <cjk>
	`桶`: [u8(0x89), 0xB1] // U+6876 <cjk>
	`牡`: [u8(0x89), 0xB2] // U+7261 <cjk>
	`乙`: [u8(0x89), 0xB3] // U+4E59 <cjk>
	`俺`: [u8(0x89), 0xB4] // U+4FFA <cjk>
	`卸`: [u8(0x89), 0xB5] // U+5378 <cjk>
	`恩`: [u8(0x89), 0xB6] // U+6069 <cjk>
	`温`: [u8(0x89), 0xB7] // U+6E29 <cjk>
	`穏`: [u8(0x89), 0xB8] // U+7A4F <cjk>
	`音`: [u8(0x89), 0xB9] // U+97F3 <cjk>
	`下`: [u8(0x89), 0xBA] // U+4E0B <cjk>
	`化`: [u8(0x89), 0xBB] // U+5316 <cjk>
	`仮`: [u8(0x89), 0xBC] // U+4EEE <cjk>
	`何`: [u8(0x89), 0xBD] // U+4F55 <cjk>
	`伽`: [u8(0x89), 0xBE] // U+4F3D <cjk>
	`価`: [u8(0x89), 0xBF] // U+4FA1 <cjk>
	`佳`: [u8(0x89), 0xC0] // U+4F73 <cjk>
	`加`: [u8(0x89), 0xC1] // U+52A0 <cjk>
	`可`: [u8(0x89), 0xC2] // U+53EF <cjk>
	`嘉`: [u8(0x89), 0xC3] // U+5609 <cjk>
	`夏`: [u8(0x89), 0xC4] // U+590F <cjk>
	`嫁`: [u8(0x89), 0xC5] // U+5AC1 <cjk>
	`家`: [u8(0x89), 0xC6] // U+5BB6 <cjk>
	`寡`: [u8(0x89), 0xC7] // U+5BE1 <cjk>
	`科`: [u8(0x89), 0xC8] // U+79D1 <cjk>
	`暇`: [u8(0x89), 0xC9] // U+6687 <cjk>
	`果`: [u8(0x89), 0xCA] // U+679C <cjk>
	`架`: [u8(0x89), 0xCB] // U+67B6 <cjk>
	`歌`: [u8(0x89), 0xCC] // U+6B4C <cjk>
	`河`: [u8(0x89), 0xCD] // U+6CB3 <cjk>
	`火`: [u8(0x89), 0xCE] // U+706B <cjk>
	`珂`: [u8(0x89), 0xCF] // U+73C2 <cjk>
	`禍`: [u8(0x89), 0xD0] // U+798D <cjk>
	`禾`: [u8(0x89), 0xD1] // U+79BE <cjk>
	`稼`: [u8(0x89), 0xD2] // U+7A3C <cjk>
	`箇`: [u8(0x89), 0xD3] // U+7B87 <cjk>
	`花`: [u8(0x89), 0xD4] // U+82B1 <cjk>
	`苛`: [u8(0x89), 0xD5] // U+82DB <cjk>
	`茄`: [u8(0x89), 0xD6] // U+8304 <cjk>
	`荷`: [u8(0x89), 0xD7] // U+8377 <cjk>
	`華`: [u8(0x89), 0xD8] // U+83EF <cjk>
	`菓`: [u8(0x89), 0xD9] // U+83D3 <cjk>
	`蝦`: [u8(0x89), 0xDA] // U+8766 <cjk>
	`課`: [u8(0x89), 0xDB] // U+8AB2 <cjk>
	`嘩`: [u8(0x89), 0xDC] // U+5629 <cjk>
	`貨`: [u8(0x89), 0xDD] // U+8CA8 <cjk>
	`迦`: [u8(0x89), 0xDE] // U+8FE6 <cjk>
	`過`: [u8(0x89), 0xDF] // U+904E <cjk>
	`霞`: [u8(0x89), 0xE0] // U+971E <cjk>
	`蚊`: [u8(0x89), 0xE1] // U+868A <cjk>
	`俄`: [u8(0x89), 0xE2] // U+4FC4 <cjk>
	`峨`: [u8(0x89), 0xE3] // U+5CE8 <cjk>
	`我`: [u8(0x89), 0xE4] // U+6211 <cjk>
	`牙`: [u8(0x89), 0xE5] // U+7259 <cjk>
	`画`: [u8(0x89), 0xE6] // U+753B <cjk>
	`臥`: [u8(0x89), 0xE7] // U+81E5 <cjk>
	`芽`: [u8(0x89), 0xE8] // U+82BD <cjk>
	`蛾`: [u8(0x89), 0xE9] // U+86FE <cjk>
	`賀`: [u8(0x89), 0xEA] // U+8CC0 <cjk>
	`雅`: [u8(0x89), 0xEB] // U+96C5 <cjk>
	`餓`: [u8(0x89), 0xEC] // U+9913 <cjk>
	`駕`: [u8(0x89), 0xED] // U+99D5 <cjk>
	`介`: [u8(0x89), 0xEE] // U+4ECB <cjk>
	`会`: [u8(0x89), 0xEF] // U+4F1A <cjk>
	`解`: [u8(0x89), 0xF0] // U+89E3 <cjk>
	`回`: [u8(0x89), 0xF1] // U+56DE <cjk>
	`塊`: [u8(0x89), 0xF2] // U+584A <cjk>
	`壊`: [u8(0x89), 0xF3] // U+58CA <cjk>
	`廻`: [u8(0x89), 0xF4] // U+5EFB <cjk>
	`快`: [u8(0x89), 0xF5] // U+5FEB <cjk>
	`怪`: [u8(0x89), 0xF6] // U+602A <cjk>
	`悔`: [u8(0x89), 0xF7] // U+6094 <cjk>
	`恢`: [u8(0x89), 0xF8] // U+6062 <cjk>
	`懐`: [u8(0x89), 0xF9] // U+61D0 <cjk>
	`戒`: [u8(0x89), 0xFA] // U+6212 <cjk>
	`拐`: [u8(0x89), 0xFB] // U+62D0 <cjk>
	`改`: [u8(0x89), 0xFC] // U+6539 <cjk>
	`魁`: [u8(0x8A), 0x40] // U+9B41 <cjk>
	`晦`: [u8(0x8A), 0x41] // U+6666 <cjk>
	`械`: [u8(0x8A), 0x42] // U+68B0 <cjk>
	`海`: [u8(0x8A), 0x43] // U+6D77 <cjk>
	`灰`: [u8(0x8A), 0x44] // U+7070 <cjk>
	`界`: [u8(0x8A), 0x45] // U+754C <cjk>
	`皆`: [u8(0x8A), 0x46] // U+7686 <cjk>
	`絵`: [u8(0x8A), 0x47] // U+7D75 <cjk>
	`芥`: [u8(0x8A), 0x48] // U+82A5 <cjk>
	`蟹`: [u8(0x8A), 0x49] // U+87F9 <cjk>
	`開`: [u8(0x8A), 0x4A] // U+958B <cjk>
	`階`: [u8(0x8A), 0x4B] // U+968E <cjk>
	`貝`: [u8(0x8A), 0x4C] // U+8C9D <cjk>
	`凱`: [u8(0x8A), 0x4D] // U+51F1 <cjk>
	`劾`: [u8(0x8A), 0x4E] // U+52BE <cjk>
	`外`: [u8(0x8A), 0x4F] // U+5916 <cjk>
	`咳`: [u8(0x8A), 0x50] // U+54B3 <cjk>
	`害`: [u8(0x8A), 0x51] // U+5BB3 <cjk>
	`崖`: [u8(0x8A), 0x52] // U+5D16 <cjk>
	`慨`: [u8(0x8A), 0x53] // U+6168 <cjk>
	`概`: [u8(0x8A), 0x54] // U+6982 <cjk>
	`涯`: [u8(0x8A), 0x55] // U+6DAF <cjk>
	`碍`: [u8(0x8A), 0x56] // U+788D <cjk>
	`蓋`: [u8(0x8A), 0x57] // U+84CB <cjk>
	`街`: [u8(0x8A), 0x58] // U+8857 <cjk>
	`該`: [u8(0x8A), 0x59] // U+8A72 <cjk>
	`鎧`: [u8(0x8A), 0x5A] // U+93A7 <cjk>
	`骸`: [u8(0x8A), 0x5B] // U+9AB8 <cjk>
	`浬`: [u8(0x8A), 0x5C] // U+6D6C <cjk>
	`馨`: [u8(0x8A), 0x5D] // U+99A8 <cjk>
	`蛙`: [u8(0x8A), 0x5E] // U+86D9 <cjk>
	`垣`: [u8(0x8A), 0x5F] // U+57A3 <cjk>
	`柿`: [u8(0x8A), 0x60] // U+67FF <cjk>
	`蛎`: [u8(0x8A), 0x61] // U+86CE <cjk>
	`鈎`: [u8(0x8A), 0x62] // U+920E <cjk>
	`劃`: [u8(0x8A), 0x63] // U+5283 <cjk>
	`嚇`: [u8(0x8A), 0x64] // U+5687 <cjk>
	`各`: [u8(0x8A), 0x65] // U+5404 <cjk>
	`廓`: [u8(0x8A), 0x66] // U+5ED3 <cjk>
	`拡`: [u8(0x8A), 0x67] // U+62E1 <cjk>
	`撹`: [u8(0x8A), 0x68] // U+64B9 <cjk>
	`格`: [u8(0x8A), 0x69] // U+683C <cjk>
	`核`: [u8(0x8A), 0x6A] // U+6838 <cjk>
	`殻`: [u8(0x8A), 0x6B] // U+6BBB <cjk>
	`獲`: [u8(0x8A), 0x6C] // U+7372 <cjk>
	`確`: [u8(0x8A), 0x6D] // U+78BA <cjk>
	`穫`: [u8(0x8A), 0x6E] // U+7A6B <cjk>
	`覚`: [u8(0x8A), 0x6F] // U+899A <cjk>
	`角`: [u8(0x8A), 0x70] // U+89D2 <cjk>
	`赫`: [u8(0x8A), 0x71] // U+8D6B <cjk>
	`較`: [u8(0x8A), 0x72] // U+8F03 <cjk>
	`郭`: [u8(0x8A), 0x73] // U+90ED <cjk>
	`閣`: [u8(0x8A), 0x74] // U+95A3 <cjk>
	`隔`: [u8(0x8A), 0x75] // U+9694 <cjk>
	`革`: [u8(0x8A), 0x76] // U+9769 <cjk>
	`学`: [u8(0x8A), 0x77] // U+5B66 <cjk>
	`岳`: [u8(0x8A), 0x78] // U+5CB3 <cjk>
	`楽`: [u8(0x8A), 0x79] // U+697D <cjk>
	`額`: [u8(0x8A), 0x7A] // U+984D <cjk>
	`顎`: [u8(0x8A), 0x7B] // U+984E <cjk>
	`掛`: [u8(0x8A), 0x7C] // U+639B <cjk>
	`笠`: [u8(0x8A), 0x7D] // U+7B20 <cjk>
	`樫`: [u8(0x8A), 0x7E] // U+6A2B <cjk>
	`橿`: [u8(0x8A), 0x80] // U+6A7F <cjk>
	`梶`: [u8(0x8A), 0x81] // U+68B6 <cjk>
	`鰍`: [u8(0x8A), 0x82] // U+9C0D <cjk>
	`潟`: [u8(0x8A), 0x83] // U+6F5F <cjk>
	`割`: [u8(0x8A), 0x84] // U+5272 <cjk>
	`喝`: [u8(0x8A), 0x85] // U+559D <cjk>
	`恰`: [u8(0x8A), 0x86] // U+6070 <cjk>
	`括`: [u8(0x8A), 0x87] // U+62EC <cjk>
	`活`: [u8(0x8A), 0x88] // U+6D3B <cjk>
	`渇`: [u8(0x8A), 0x89] // U+6E07 <cjk>
	`滑`: [u8(0x8A), 0x8A] // U+6ED1 <cjk>
	`葛`: [u8(0x8A), 0x8B] // U+845B <cjk>
	`褐`: [u8(0x8A), 0x8C] // U+8910 <cjk>
	`轄`: [u8(0x8A), 0x8D] // U+8F44 <cjk>
	`且`: [u8(0x8A), 0x8E] // U+4E14 <cjk>
	`鰹`: [u8(0x8A), 0x8F] // U+9C39 <cjk>
	`叶`: [u8(0x8A), 0x90] // U+53F6 <cjk>
	`椛`: [u8(0x8A), 0x91] // U+691B <cjk>
	`樺`: [u8(0x8A), 0x92] // U+6A3A <cjk>
	`鞄`: [u8(0x8A), 0x93] // U+9784 <cjk>
	`株`: [u8(0x8A), 0x94] // U+682A <cjk>
	`兜`: [u8(0x8A), 0x95] // U+515C <cjk>
	`竃`: [u8(0x8A), 0x96] // U+7AC3 <cjk>
	`蒲`: [u8(0x8A), 0x97] // U+84B2 <cjk>
	`釜`: [u8(0x8A), 0x98] // U+91DC <cjk>
	`鎌`: [u8(0x8A), 0x99] // U+938C <cjk>
	`噛`: [u8(0x8A), 0x9A] // U+565B <cjk>
	`鴨`: [u8(0x8A), 0x9B] // U+9D28 <cjk>
	`栢`: [u8(0x8A), 0x9C] // U+6822 <cjk>
	`茅`: [u8(0x8A), 0x9D] // U+8305 <cjk>
	`萱`: [u8(0x8A), 0x9E] // U+8431 <cjk>
	`粥`: [u8(0x8A), 0x9F] // U+7CA5 <cjk>
	`刈`: [u8(0x8A), 0xA0] // U+5208 <cjk>
	`苅`: [u8(0x8A), 0xA1] // U+82C5 <cjk>
	`瓦`: [u8(0x8A), 0xA2] // U+74E6 <cjk>
	`乾`: [u8(0x8A), 0xA3] // U+4E7E <cjk>
	`侃`: [u8(0x8A), 0xA4] // U+4F83 <cjk>
	`冠`: [u8(0x8A), 0xA5] // U+51A0 <cjk>
	`寒`: [u8(0x8A), 0xA6] // U+5BD2 <cjk>
	`刊`: [u8(0x8A), 0xA7] // U+520A <cjk>
	`勘`: [u8(0x8A), 0xA8] // U+52D8 <cjk>
	`勧`: [u8(0x8A), 0xA9] // U+52E7 <cjk>
	`巻`: [u8(0x8A), 0xAA] // U+5DFB <cjk>
	`喚`: [u8(0x8A), 0xAB] // U+559A <cjk>
	`堪`: [u8(0x8A), 0xAC] // U+582A <cjk>
	`姦`: [u8(0x8A), 0xAD] // U+59E6 <cjk>
	`完`: [u8(0x8A), 0xAE] // U+5B8C <cjk>
	`官`: [u8(0x8A), 0xAF] // U+5B98 <cjk>
	`寛`: [u8(0x8A), 0xB0] // U+5BDB <cjk>
	`干`: [u8(0x8A), 0xB1] // U+5E72 <cjk>
	`幹`: [u8(0x8A), 0xB2] // U+5E79 <cjk>
	`患`: [u8(0x8A), 0xB3] // U+60A3 <cjk>
	`感`: [u8(0x8A), 0xB4] // U+611F <cjk>
	`慣`: [u8(0x8A), 0xB5] // U+6163 <cjk>
	`憾`: [u8(0x8A), 0xB6] // U+61BE <cjk>
	`換`: [u8(0x8A), 0xB7] // U+63DB <cjk>
	`敢`: [u8(0x8A), 0xB8] // U+6562 <cjk>
	`柑`: [u8(0x8A), 0xB9] // U+67D1 <cjk>
	`桓`: [u8(0x8A), 0xBA] // U+6853 <cjk>
	`棺`: [u8(0x8A), 0xBB] // U+68FA <cjk>
	`款`: [u8(0x8A), 0xBC] // U+6B3E <cjk>
	`歓`: [u8(0x8A), 0xBD] // U+6B53 <cjk>
	`汗`: [u8(0x8A), 0xBE] // U+6C57 <cjk>
	`漢`: [u8(0x8A), 0xBF] // U+6F22 <cjk>
	`澗`: [u8(0x8A), 0xC0] // U+6F97 <cjk>
	`潅`: [u8(0x8A), 0xC1] // U+6F45 <cjk>
	`環`: [u8(0x8A), 0xC2] // U+74B0 <cjk>
	`甘`: [u8(0x8A), 0xC3] // U+7518 <cjk>
	`監`: [u8(0x8A), 0xC4] // U+76E3 <cjk>
	`看`: [u8(0x8A), 0xC5] // U+770B <cjk>
	`竿`: [u8(0x8A), 0xC6] // U+7AFF <cjk>
	`管`: [u8(0x8A), 0xC7] // U+7BA1 <cjk>
	`簡`: [u8(0x8A), 0xC8] // U+7C21 <cjk>
	`緩`: [u8(0x8A), 0xC9] // U+7DE9 <cjk>
	`缶`: [u8(0x8A), 0xCA] // U+7F36 <cjk>
	`翰`: [u8(0x8A), 0xCB] // U+7FF0 <cjk>
	`肝`: [u8(0x8A), 0xCC] // U+809D <cjk>
	`艦`: [u8(0x8A), 0xCD] // U+8266 <cjk>
	`莞`: [u8(0x8A), 0xCE] // U+839E <cjk>
	`観`: [u8(0x8A), 0xCF] // U+89B3 <cjk>
	`諌`: [u8(0x8A), 0xD0] // U+8ACC <cjk>
	`貫`: [u8(0x8A), 0xD1] // U+8CAB <cjk>
	`還`: [u8(0x8A), 0xD2] // U+9084 <cjk>
	`鑑`: [u8(0x8A), 0xD3] // U+9451 <cjk>
	`間`: [u8(0x8A), 0xD4] // U+9593 <cjk>
	`閑`: [u8(0x8A), 0xD5] // U+9591 <cjk>
	`関`: [u8(0x8A), 0xD6] // U+95A2 <cjk>
	`陥`: [u8(0x8A), 0xD7] // U+9665 <cjk>
	`韓`: [u8(0x8A), 0xD8] // U+97D3 <cjk>
	`館`: [u8(0x8A), 0xD9] // U+9928 <cjk>
	`舘`: [u8(0x8A), 0xDA] // U+8218 <cjk>
	`丸`: [u8(0x8A), 0xDB] // U+4E38 <cjk>
	`含`: [u8(0x8A), 0xDC] // U+542B <cjk>
	`岸`: [u8(0x8A), 0xDD] // U+5CB8 <cjk>
	`巌`: [u8(0x8A), 0xDE] // U+5DCC <cjk>
	`玩`: [u8(0x8A), 0xDF] // U+73A9 <cjk>
	`癌`: [u8(0x8A), 0xE0] // U+764C <cjk>
	`眼`: [u8(0x8A), 0xE1] // U+773C <cjk>
	`岩`: [u8(0x8A), 0xE2] // U+5CA9 <cjk>
	`翫`: [u8(0x8A), 0xE3] // U+7FEB <cjk>
	`贋`: [u8(0x8A), 0xE4] // U+8D0B <cjk>
	`雁`: [u8(0x8A), 0xE5] // U+96C1 <cjk>
	`頑`: [u8(0x8A), 0xE6] // U+9811 <cjk>
	`顔`: [u8(0x8A), 0xE7] // U+9854 <cjk>
	`願`: [u8(0x8A), 0xE8] // U+9858 <cjk>
	`企`: [u8(0x8A), 0xE9] // U+4F01 <cjk>
	`伎`: [u8(0x8A), 0xEA] // U+4F0E <cjk>
	`危`: [u8(0x8A), 0xEB] // U+5371 <cjk>
	`喜`: [u8(0x8A), 0xEC] // U+559C <cjk>
	`器`: [u8(0x8A), 0xED] // U+5668 <cjk>
	`基`: [u8(0x8A), 0xEE] // U+57FA <cjk>
	`奇`: [u8(0x8A), 0xEF] // U+5947 <cjk>
	`嬉`: [u8(0x8A), 0xF0] // U+5B09 <cjk>
	`寄`: [u8(0x8A), 0xF1] // U+5BC4 <cjk>
	`岐`: [u8(0x8A), 0xF2] // U+5C90 <cjk>
	`希`: [u8(0x8A), 0xF3] // U+5E0C <cjk>
	`幾`: [u8(0x8A), 0xF4] // U+5E7E <cjk>
	`忌`: [u8(0x8A), 0xF5] // U+5FCC <cjk>
	`揮`: [u8(0x8A), 0xF6] // U+63EE <cjk>
	`机`: [u8(0x8A), 0xF7] // U+673A <cjk>
	`旗`: [u8(0x8A), 0xF8] // U+65D7 <cjk>
	`既`: [u8(0x8A), 0xF9] // U+65E2 <cjk>
	`期`: [u8(0x8A), 0xFA] // U+671F <cjk>
	`棋`: [u8(0x8A), 0xFB] // U+68CB <cjk>
	`棄`: [u8(0x8A), 0xFC] // U+68C4 <cjk>
	`機`: [u8(0x8B), 0x40] // U+6A5F <cjk>
	`帰`: [u8(0x8B), 0x41] // U+5E30 <cjk>
	`毅`: [u8(0x8B), 0x42] // U+6BC5 <cjk>
	`気`: [u8(0x8B), 0x43] // U+6C17 <cjk>
	`汽`: [u8(0x8B), 0x44] // U+6C7D <cjk>
	`畿`: [u8(0x8B), 0x45] // U+757F <cjk>
	`祈`: [u8(0x8B), 0x46] // U+7948 <cjk>
	`季`: [u8(0x8B), 0x47] // U+5B63 <cjk>
	`稀`: [u8(0x8B), 0x48] // U+7A00 <cjk>
	`紀`: [u8(0x8B), 0x49] // U+7D00 <cjk>
	`徽`: [u8(0x8B), 0x4A] // U+5FBD <cjk>
	`規`: [u8(0x8B), 0x4B] // U+898F <cjk>
	`記`: [u8(0x8B), 0x4C] // U+8A18 <cjk>
	`貴`: [u8(0x8B), 0x4D] // U+8CB4 <cjk>
	`起`: [u8(0x8B), 0x4E] // U+8D77 <cjk>
	`軌`: [u8(0x8B), 0x4F] // U+8ECC <cjk>
	`輝`: [u8(0x8B), 0x50] // U+8F1D <cjk>
	`飢`: [u8(0x8B), 0x51] // U+98E2 <cjk>
	`騎`: [u8(0x8B), 0x52] // U+9A0E <cjk>
	`鬼`: [u8(0x8B), 0x53] // U+9B3C <cjk>
	`亀`: [u8(0x8B), 0x54] // U+4E80 <cjk>
	`偽`: [u8(0x8B), 0x55] // U+507D <cjk>
	`儀`: [u8(0x8B), 0x56] // U+5100 <cjk>
	`妓`: [u8(0x8B), 0x57] // U+5993 <cjk>
	`宜`: [u8(0x8B), 0x58] // U+5B9C <cjk>
	`戯`: [u8(0x8B), 0x59] // U+622F <cjk>
	`技`: [u8(0x8B), 0x5A] // U+6280 <cjk>
	`擬`: [u8(0x8B), 0x5B] // U+64EC <cjk>
	`欺`: [u8(0x8B), 0x5C] // U+6B3A <cjk>
	`犠`: [u8(0x8B), 0x5D] // U+72A0 <cjk>
	`疑`: [u8(0x8B), 0x5E] // U+7591 <cjk>
	`祇`: [u8(0x8B), 0x5F] // U+7947 <cjk>
	`義`: [u8(0x8B), 0x60] // U+7FA9 <cjk>
	`蟻`: [u8(0x8B), 0x61] // U+87FB <cjk>
	`誼`: [u8(0x8B), 0x62] // U+8ABC <cjk>
	`議`: [u8(0x8B), 0x63] // U+8B70 <cjk>
	`掬`: [u8(0x8B), 0x64] // U+63AC <cjk>
	`菊`: [u8(0x8B), 0x65] // U+83CA <cjk>
	`鞠`: [u8(0x8B), 0x66] // U+97A0 <cjk>
	`吉`: [u8(0x8B), 0x67] // U+5409 <cjk>
	`吃`: [u8(0x8B), 0x68] // U+5403 <cjk>
	`喫`: [u8(0x8B), 0x69] // U+55AB <cjk>
	`桔`: [u8(0x8B), 0x6A] // U+6854 <cjk>
	`橘`: [u8(0x8B), 0x6B] // U+6A58 <cjk>
	`詰`: [u8(0x8B), 0x6C] // U+8A70 <cjk>
	`砧`: [u8(0x8B), 0x6D] // U+7827 <cjk>
	`杵`: [u8(0x8B), 0x6E] // U+6775 <cjk>
	`黍`: [u8(0x8B), 0x6F] // U+9ECD <cjk>
	`却`: [u8(0x8B), 0x70] // U+5374 <cjk>
	`客`: [u8(0x8B), 0x71] // U+5BA2 <cjk>
	`脚`: [u8(0x8B), 0x72] // U+811A <cjk>
	`虐`: [u8(0x8B), 0x73] // U+8650 <cjk>
	`逆`: [u8(0x8B), 0x74] // U+9006 <cjk>
	`丘`: [u8(0x8B), 0x75] // U+4E18 <cjk>
	`久`: [u8(0x8B), 0x76] // U+4E45 <cjk>
	`仇`: [u8(0x8B), 0x77] // U+4EC7 <cjk>
	`休`: [u8(0x8B), 0x78] // U+4F11 <cjk>
	`及`: [u8(0x8B), 0x79] // U+53CA <cjk>
	`吸`: [u8(0x8B), 0x7A] // U+5438 <cjk>
	`宮`: [u8(0x8B), 0x7B] // U+5BAE <cjk>
	`弓`: [u8(0x8B), 0x7C] // U+5F13 <cjk>
	`急`: [u8(0x8B), 0x7D] // U+6025 <cjk>
	`救`: [u8(0x8B), 0x7E] // U+6551 <cjk>
	`朽`: [u8(0x8B), 0x80] // U+673D <cjk>
	`求`: [u8(0x8B), 0x81] // U+6C42 <cjk>
	`汲`: [u8(0x8B), 0x82] // U+6C72 <cjk>
	`泣`: [u8(0x8B), 0x83] // U+6CE3 <cjk>
	`灸`: [u8(0x8B), 0x84] // U+7078 <cjk>
	`球`: [u8(0x8B), 0x85] // U+7403 <cjk>
	`究`: [u8(0x8B), 0x86] // U+7A76 <cjk>
	`窮`: [u8(0x8B), 0x87] // U+7AAE <cjk>
	`笈`: [u8(0x8B), 0x88] // U+7B08 <cjk>
	`級`: [u8(0x8B), 0x89] // U+7D1A <cjk>
	`糾`: [u8(0x8B), 0x8A] // U+7CFE <cjk>
	`給`: [u8(0x8B), 0x8B] // U+7D66 <cjk>
	`旧`: [u8(0x8B), 0x8C] // U+65E7 <cjk>
	`牛`: [u8(0x8B), 0x8D] // U+725B <cjk>
	`去`: [u8(0x8B), 0x8E] // U+53BB <cjk>
	`居`: [u8(0x8B), 0x8F] // U+5C45 <cjk>
	`巨`: [u8(0x8B), 0x90] // U+5DE8 <cjk>
	`拒`: [u8(0x8B), 0x91] // U+62D2 <cjk>
	`拠`: [u8(0x8B), 0x92] // U+62E0 <cjk>
	`挙`: [u8(0x8B), 0x93] // U+6319 <cjk>
	`渠`: [u8(0x8B), 0x94] // U+6E20 <cjk>
	`虚`: [u8(0x8B), 0x95] // U+865A <cjk>
	`許`: [u8(0x8B), 0x96] // U+8A31 <cjk>
	`距`: [u8(0x8B), 0x97] // U+8DDD <cjk>
	`鋸`: [u8(0x8B), 0x98] // U+92F8 <cjk>
	`漁`: [u8(0x8B), 0x99] // U+6F01 <cjk>
	`禦`: [u8(0x8B), 0x9A] // U+79A6 <cjk>
	`魚`: [u8(0x8B), 0x9B] // U+9B5A <cjk>
	`亨`: [u8(0x8B), 0x9C] // U+4EA8 <cjk>
	`享`: [u8(0x8B), 0x9D] // U+4EAB <cjk>
	`京`: [u8(0x8B), 0x9E] // U+4EAC <cjk>
	`供`: [u8(0x8B), 0x9F] // U+4F9B <cjk>
	`侠`: [u8(0x8B), 0xA0] // U+4FA0 <cjk>
	`僑`: [u8(0x8B), 0xA1] // U+50D1 <cjk>
	`兇`: [u8(0x8B), 0xA2] // U+5147 <cjk>
	`競`: [u8(0x8B), 0xA3] // U+7AF6 <cjk>
	`共`: [u8(0x8B), 0xA4] // U+5171 <cjk>
	`凶`: [u8(0x8B), 0xA5] // U+51F6 <cjk>
	`協`: [u8(0x8B), 0xA6] // U+5354 <cjk>
	`匡`: [u8(0x8B), 0xA7] // U+5321 <cjk>
	`卿`: [u8(0x8B), 0xA8] // U+537F <cjk>
	`叫`: [u8(0x8B), 0xA9] // U+53EB <cjk>
	`喬`: [u8(0x8B), 0xAA] // U+55AC <cjk>
	`境`: [u8(0x8B), 0xAB] // U+5883 <cjk>
	`峡`: [u8(0x8B), 0xAC] // U+5CE1 <cjk>
	`強`: [u8(0x8B), 0xAD] // U+5F37 <cjk>
	`彊`: [u8(0x8B), 0xAE] // U+5F4A <cjk>
	`怯`: [u8(0x8B), 0xAF] // U+602F <cjk>
	`恐`: [u8(0x8B), 0xB0] // U+6050 <cjk>
	`恭`: [u8(0x8B), 0xB1] // U+606D <cjk>
	`挟`: [u8(0x8B), 0xB2] // U+631F <cjk>
	`教`: [u8(0x8B), 0xB3] // U+6559 <cjk>
	`橋`: [u8(0x8B), 0xB4] // U+6A4B <cjk>
	`況`: [u8(0x8B), 0xB5] // U+6CC1 <cjk>
	`狂`: [u8(0x8B), 0xB6] // U+72C2 <cjk>
	`狭`: [u8(0x8B), 0xB7] // U+72ED <cjk>
	`矯`: [u8(0x8B), 0xB8] // U+77EF <cjk>
	`胸`: [u8(0x8B), 0xB9] // U+80F8 <cjk>
	`脅`: [u8(0x8B), 0xBA] // U+8105 <cjk>
	`興`: [u8(0x8B), 0xBB] // U+8208 <cjk>
	`蕎`: [u8(0x8B), 0xBC] // U+854E <cjk>
	`郷`: [u8(0x8B), 0xBD] // U+90F7 <cjk>
	`鏡`: [u8(0x8B), 0xBE] // U+93E1 <cjk>
	`響`: [u8(0x8B), 0xBF] // U+97FF <cjk>
	`饗`: [u8(0x8B), 0xC0] // U+9957 <cjk>
	`驚`: [u8(0x8B), 0xC1] // U+9A5A <cjk>
	`仰`: [u8(0x8B), 0xC2] // U+4EF0 <cjk>
	`凝`: [u8(0x8B), 0xC3] // U+51DD <cjk>
	`尭`: [u8(0x8B), 0xC4] // U+5C2D <cjk>
	`暁`: [u8(0x8B), 0xC5] // U+6681 <cjk>
	`業`: [u8(0x8B), 0xC6] // U+696D <cjk>
	`局`: [u8(0x8B), 0xC7] // U+5C40 <cjk>
	`曲`: [u8(0x8B), 0xC8] // U+66F2 <cjk>
	`極`: [u8(0x8B), 0xC9] // U+6975 <cjk>
	`玉`: [u8(0x8B), 0xCA] // U+7389 <cjk>
	`桐`: [u8(0x8B), 0xCB] // U+6850 <cjk>
	`粁`: [u8(0x8B), 0xCC] // U+7C81 <cjk>
	`僅`: [u8(0x8B), 0xCD] // U+50C5 <cjk>
	`勤`: [u8(0x8B), 0xCE] // U+52E4 <cjk>
	`均`: [u8(0x8B), 0xCF] // U+5747 <cjk>
	`巾`: [u8(0x8B), 0xD0] // U+5DFE <cjk>
	`錦`: [u8(0x8B), 0xD1] // U+9326 <cjk>
	`斤`: [u8(0x8B), 0xD2] // U+65A4 <cjk>
	`欣`: [u8(0x8B), 0xD3] // U+6B23 <cjk>
	`欽`: [u8(0x8B), 0xD4] // U+6B3D <cjk>
	`琴`: [u8(0x8B), 0xD5] // U+7434 <cjk>
	`禁`: [u8(0x8B), 0xD6] // U+7981 <cjk>
	`禽`: [u8(0x8B), 0xD7] // U+79BD <cjk>
	`筋`: [u8(0x8B), 0xD8] // U+7B4B <cjk>
	`緊`: [u8(0x8B), 0xD9] // U+7DCA <cjk>
	`芹`: [u8(0x8B), 0xDA] // U+82B9 <cjk>
	`菌`: [u8(0x8B), 0xDB] // U+83CC <cjk>
	`衿`: [u8(0x8B), 0xDC] // U+887F <cjk>
	`襟`: [u8(0x8B), 0xDD] // U+895F <cjk>
	`謹`: [u8(0x8B), 0xDE] // U+8B39 <cjk>
	`近`: [u8(0x8B), 0xDF] // U+8FD1 <cjk>
	`金`: [u8(0x8B), 0xE0] // U+91D1 <cjk>
	`吟`: [u8(0x8B), 0xE1] // U+541F <cjk>
	`銀`: [u8(0x8B), 0xE2] // U+9280 <cjk>
	`九`: [u8(0x8B), 0xE3] // U+4E5D <cjk>
	`倶`: [u8(0x8B), 0xE4] // U+5036 <cjk>
	`句`: [u8(0x8B), 0xE5] // U+53E5 <cjk>
	`区`: [u8(0x8B), 0xE6] // U+533A <cjk>
	`狗`: [u8(0x8B), 0xE7] // U+72D7 <cjk>
	`玖`: [u8(0x8B), 0xE8] // U+7396 <cjk>
	`矩`: [u8(0x8B), 0xE9] // U+77E9 <cjk>
	`苦`: [u8(0x8B), 0xEA] // U+82E6 <cjk>
	`躯`: [u8(0x8B), 0xEB] // U+8EAF <cjk>
	`駆`: [u8(0x8B), 0xEC] // U+99C6 <cjk>
	`駈`: [u8(0x8B), 0xED] // U+99C8 <cjk>
	`駒`: [u8(0x8B), 0xEE] // U+99D2 <cjk>
	`具`: [u8(0x8B), 0xEF] // U+5177 <cjk>
	`愚`: [u8(0x8B), 0xF0] // U+611A <cjk>
	`虞`: [u8(0x8B), 0xF1] // U+865E <cjk>
	`喰`: [u8(0x8B), 0xF2] // U+55B0 <cjk>
	`空`: [u8(0x8B), 0xF3] // U+7A7A <cjk>
	`偶`: [u8(0x8B), 0xF4] // U+5076 <cjk>
	`寓`: [u8(0x8B), 0xF5] // U+5BD3 <cjk>
	`遇`: [u8(0x8B), 0xF6] // U+9047 <cjk>
	`隅`: [u8(0x8B), 0xF7] // U+9685 <cjk>
	`串`: [u8(0x8B), 0xF8] // U+4E32 <cjk>
	`櫛`: [u8(0x8B), 0xF9] // U+6ADB <cjk>
	`釧`: [u8(0x8B), 0xFA] // U+91E7 <cjk>
	`屑`: [u8(0x8B), 0xFB] // U+5C51 <cjk>
	`屈`: [u8(0x8B), 0xFC] // U+5C48 <cjk>
	`掘`: [u8(0x8C), 0x40] // U+6398 <cjk>
	`窟`: [u8(0x8C), 0x41] // U+7A9F <cjk>
	`沓`: [u8(0x8C), 0x42] // U+6C93 <cjk>
	`靴`: [u8(0x8C), 0x43] // U+9774 <cjk>
	`轡`: [u8(0x8C), 0x44] // U+8F61 <cjk>
	`窪`: [u8(0x8C), 0x45] // U+7AAA <cjk>
	`熊`: [u8(0x8C), 0x46] // U+718A <cjk>
	`隈`: [u8(0x8C), 0x47] // U+9688 <cjk>
	`粂`: [u8(0x8C), 0x48] // U+7C82 <cjk>
	`栗`: [u8(0x8C), 0x49] // U+6817 <cjk>
	`繰`: [u8(0x8C), 0x4A] // U+7E70 <cjk>
	`桑`: [u8(0x8C), 0x4B] // U+6851 <cjk>
	`鍬`: [u8(0x8C), 0x4C] // U+936C <cjk>
	`勲`: [u8(0x8C), 0x4D] // U+52F2 <cjk>
	`君`: [u8(0x8C), 0x4E] // U+541B <cjk>
	`薫`: [u8(0x8C), 0x4F] // U+85AB <cjk>
	`訓`: [u8(0x8C), 0x50] // U+8A13 <cjk>
	`群`: [u8(0x8C), 0x51] // U+7FA4 <cjk>
	`軍`: [u8(0x8C), 0x52] // U+8ECD <cjk>
	`郡`: [u8(0x8C), 0x53] // U+90E1 <cjk>
	`卦`: [u8(0x8C), 0x54] // U+5366 <cjk>
	`袈`: [u8(0x8C), 0x55] // U+8888 <cjk>
	`祁`: [u8(0x8C), 0x56] // U+7941 <cjk>
	`係`: [u8(0x8C), 0x57] // U+4FC2 <cjk>
	`傾`: [u8(0x8C), 0x58] // U+50BE <cjk>
	`刑`: [u8(0x8C), 0x59] // U+5211 <cjk>
	`兄`: [u8(0x8C), 0x5A] // U+5144 <cjk>
	`啓`: [u8(0x8C), 0x5B] // U+5553 <cjk>
	`圭`: [u8(0x8C), 0x5C] // U+572D <cjk>
	`珪`: [u8(0x8C), 0x5D] // U+73EA <cjk>
	`型`: [u8(0x8C), 0x5E] // U+578B <cjk>
	`契`: [u8(0x8C), 0x5F] // U+5951 <cjk>
	`形`: [u8(0x8C), 0x60] // U+5F62 <cjk>
	`径`: [u8(0x8C), 0x61] // U+5F84 <cjk>
	`恵`: [u8(0x8C), 0x62] // U+6075 <cjk>
	`慶`: [u8(0x8C), 0x63] // U+6176 <cjk>
	`慧`: [u8(0x8C), 0x64] // U+6167 <cjk>
	`憩`: [u8(0x8C), 0x65] // U+61A9 <cjk>
	`掲`: [u8(0x8C), 0x66] // U+63B2 <cjk>
	`携`: [u8(0x8C), 0x67] // U+643A <cjk>
	`敬`: [u8(0x8C), 0x68] // U+656C <cjk>
	`景`: [u8(0x8C), 0x69] // U+666F <cjk>
	`桂`: [u8(0x8C), 0x6A] // U+6842 <cjk>
	`渓`: [u8(0x8C), 0x6B] // U+6E13 <cjk>
	`畦`: [u8(0x8C), 0x6C] // U+7566 <cjk>
	`稽`: [u8(0x8C), 0x6D] // U+7A3D <cjk>
	`系`: [u8(0x8C), 0x6E] // U+7CFB <cjk>
	`経`: [u8(0x8C), 0x6F] // U+7D4C <cjk>
	`継`: [u8(0x8C), 0x70] // U+7D99 <cjk>
	`繋`: [u8(0x8C), 0x71] // U+7E4B <cjk>
	`罫`: [u8(0x8C), 0x72] // U+7F6B <cjk>
	`茎`: [u8(0x8C), 0x73] // U+830E <cjk>
	`荊`: [u8(0x8C), 0x74] // U+834A <cjk>
	`蛍`: [u8(0x8C), 0x75] // U+86CD <cjk>
	`計`: [u8(0x8C), 0x76] // U+8A08 <cjk>
	`詣`: [u8(0x8C), 0x77] // U+8A63 <cjk>
	`警`: [u8(0x8C), 0x78] // U+8B66 <cjk>
	`軽`: [u8(0x8C), 0x79] // U+8EFD <cjk>
	`頚`: [u8(0x8C), 0x7A] // U+981A <cjk>
	`鶏`: [u8(0x8C), 0x7B] // U+9D8F <cjk>
	`芸`: [u8(0x8C), 0x7C] // U+82B8 <cjk>
	`迎`: [u8(0x8C), 0x7D] // U+8FCE <cjk>
	`鯨`: [u8(0x8C), 0x7E] // U+9BE8 <cjk>
	`劇`: [u8(0x8C), 0x80] // U+5287 <cjk>
	`戟`: [u8(0x8C), 0x81] // U+621F <cjk>
	`撃`: [u8(0x8C), 0x82] // U+6483 <cjk>
	`激`: [u8(0x8C), 0x83] // U+6FC0 <cjk>
	`隙`: [u8(0x8C), 0x84] // U+9699 <cjk>
	`桁`: [u8(0x8C), 0x85] // U+6841 <cjk>
	`傑`: [u8(0x8C), 0x86] // U+5091 <cjk>
	`欠`: [u8(0x8C), 0x87] // U+6B20 <cjk>
	`決`: [u8(0x8C), 0x88] // U+6C7A <cjk>
	`潔`: [u8(0x8C), 0x89] // U+6F54 <cjk>
	`穴`: [u8(0x8C), 0x8A] // U+7A74 <cjk>
	`結`: [u8(0x8C), 0x8B] // U+7D50 <cjk>
	`血`: [u8(0x8C), 0x8C] // U+8840 <cjk>
	`訣`: [u8(0x8C), 0x8D] // U+8A23 <cjk>
	`月`: [u8(0x8C), 0x8E] // U+6708 <cjk>
	`件`: [u8(0x8C), 0x8F] // U+4EF6 <cjk>
	`倹`: [u8(0x8C), 0x90] // U+5039 <cjk>
	`倦`: [u8(0x8C), 0x91] // U+5026 <cjk>
	`健`: [u8(0x8C), 0x92] // U+5065 <cjk>
	`兼`: [u8(0x8C), 0x93] // U+517C <cjk>
	`券`: [u8(0x8C), 0x94] // U+5238 <cjk>
	`剣`: [u8(0x8C), 0x95] // U+5263 <cjk>
	`喧`: [u8(0x8C), 0x96] // U+55A7 <cjk>
	`圏`: [u8(0x8C), 0x97] // U+570F <cjk>
	`堅`: [u8(0x8C), 0x98] // U+5805 <cjk>
	`嫌`: [u8(0x8C), 0x99] // U+5ACC <cjk>
	`建`: [u8(0x8C), 0x9A] // U+5EFA <cjk>
	`憲`: [u8(0x8C), 0x9B] // U+61B2 <cjk>
	`懸`: [u8(0x8C), 0x9C] // U+61F8 <cjk>
	`拳`: [u8(0x8C), 0x9D] // U+62F3 <cjk>
	`捲`: [u8(0x8C), 0x9E] // U+6372 <cjk>
	`検`: [u8(0x8C), 0x9F] // U+691C <cjk>
	`権`: [u8(0x8C), 0xA0] // U+6A29 <cjk>
	`牽`: [u8(0x8C), 0xA1] // U+727D <cjk>
	`犬`: [u8(0x8C), 0xA2] // U+72AC <cjk>
	`献`: [u8(0x8C), 0xA3] // U+732E <cjk>
	`研`: [u8(0x8C), 0xA4] // U+7814 <cjk>
	`硯`: [u8(0x8C), 0xA5] // U+786F <cjk>
	`絹`: [u8(0x8C), 0xA6] // U+7D79 <cjk>
	`県`: [u8(0x8C), 0xA7] // U+770C <cjk>
	`肩`: [u8(0x8C), 0xA8] // U+80A9 <cjk>
	`見`: [u8(0x8C), 0xA9] // U+898B <cjk>
	`謙`: [u8(0x8C), 0xAA] // U+8B19 <cjk>
	`賢`: [u8(0x8C), 0xAB] // U+8CE2 <cjk>
	`軒`: [u8(0x8C), 0xAC] // U+8ED2 <cjk>
	`遣`: [u8(0x8C), 0xAD] // U+9063 <cjk>
	`鍵`: [u8(0x8C), 0xAE] // U+9375 <cjk>
	`険`: [u8(0x8C), 0xAF] // U+967A <cjk>
	`顕`: [u8(0x8C), 0xB0] // U+9855 <cjk>
	`験`: [u8(0x8C), 0xB1] // U+9A13 <cjk>
	`鹸`: [u8(0x8C), 0xB2] // U+9E78 <cjk>
	`元`: [u8(0x8C), 0xB3] // U+5143 <cjk>
	`原`: [u8(0x8C), 0xB4] // U+539F <cjk>
	`厳`: [u8(0x8C), 0xB5] // U+53B3 <cjk>
	`幻`: [u8(0x8C), 0xB6] // U+5E7B <cjk>
	`弦`: [u8(0x8C), 0xB7] // U+5F26 <cjk>
	`減`: [u8(0x8C), 0xB8] // U+6E1B <cjk>
	`源`: [u8(0x8C), 0xB9] // U+6E90 <cjk>
	`玄`: [u8(0x8C), 0xBA] // U+7384 <cjk>
	`現`: [u8(0x8C), 0xBB] // U+73FE <cjk>
	`絃`: [u8(0x8C), 0xBC] // U+7D43 <cjk>
	`舷`: [u8(0x8C), 0xBD] // U+8237 <cjk>
	`言`: [u8(0x8C), 0xBE] // U+8A00 <cjk>
	`諺`: [u8(0x8C), 0xBF] // U+8AFA <cjk>
	`限`: [u8(0x8C), 0xC0] // U+9650 <cjk>
	`乎`: [u8(0x8C), 0xC1] // U+4E4E <cjk>
	`個`: [u8(0x8C), 0xC2] // U+500B <cjk>
	`古`: [u8(0x8C), 0xC3] // U+53E4 <cjk>
	`呼`: [u8(0x8C), 0xC4] // U+547C <cjk>
	`固`: [u8(0x8C), 0xC5] // U+56FA <cjk>
	`姑`: [u8(0x8C), 0xC6] // U+59D1 <cjk>
	`孤`: [u8(0x8C), 0xC7] // U+5B64 <cjk>
	`己`: [u8(0x8C), 0xC8] // U+5DF1 <cjk>
	`庫`: [u8(0x8C), 0xC9] // U+5EAB <cjk>
	`弧`: [u8(0x8C), 0xCA] // U+5F27 <cjk>
	`戸`: [u8(0x8C), 0xCB] // U+6238 <cjk>
	`故`: [u8(0x8C), 0xCC] // U+6545 <cjk>
	`枯`: [u8(0x8C), 0xCD] // U+67AF <cjk>
	`湖`: [u8(0x8C), 0xCE] // U+6E56 <cjk>
	`狐`: [u8(0x8C), 0xCF] // U+72D0 <cjk>
	`糊`: [u8(0x8C), 0xD0] // U+7CCA <cjk>
	`袴`: [u8(0x8C), 0xD1] // U+88B4 <cjk>
	`股`: [u8(0x8C), 0xD2] // U+80A1 <cjk>
	`胡`: [u8(0x8C), 0xD3] // U+80E1 <cjk>
	`菰`: [u8(0x8C), 0xD4] // U+83F0 <cjk>
	`虎`: [u8(0x8C), 0xD5] // U+864E <cjk>
	`誇`: [u8(0x8C), 0xD6] // U+8A87 <cjk>
	`跨`: [u8(0x8C), 0xD7] // U+8DE8 <cjk>
	`鈷`: [u8(0x8C), 0xD8] // U+9237 <cjk>
	`雇`: [u8(0x8C), 0xD9] // U+96C7 <cjk>
	`顧`: [u8(0x8C), 0xDA] // U+9867 <cjk>
	`鼓`: [u8(0x8C), 0xDB] // U+9F13 <cjk>
	`五`: [u8(0x8C), 0xDC] // U+4E94 <cjk>
	`互`: [u8(0x8C), 0xDD] // U+4E92 <cjk>
	`伍`: [u8(0x8C), 0xDE] // U+4F0D <cjk>
	`午`: [u8(0x8C), 0xDF] // U+5348 <cjk>
	`呉`: [u8(0x8C), 0xE0] // U+5449 <cjk>
	`吾`: [u8(0x8C), 0xE1] // U+543E <cjk>
	`娯`: [u8(0x8C), 0xE2] // U+5A2F <cjk>
	`後`: [u8(0x8C), 0xE3] // U+5F8C <cjk>
	`御`: [u8(0x8C), 0xE4] // U+5FA1 <cjk>
	`悟`: [u8(0x8C), 0xE5] // U+609F <cjk>
	`梧`: [u8(0x8C), 0xE6] // U+68A7 <cjk>
	`檎`: [u8(0x8C), 0xE7] // U+6A8E <cjk>
	`瑚`: [u8(0x8C), 0xE8] // U+745A <cjk>
	`碁`: [u8(0x8C), 0xE9] // U+7881 <cjk>
	`語`: [u8(0x8C), 0xEA] // U+8A9E <cjk>
	`誤`: [u8(0x8C), 0xEB] // U+8AA4 <cjk>
	`護`: [u8(0x8C), 0xEC] // U+8B77 <cjk>
	`醐`: [u8(0x8C), 0xED] // U+9190 <cjk>
	`乞`: [u8(0x8C), 0xEE] // U+4E5E <cjk>
	`鯉`: [u8(0x8C), 0xEF] // U+9BC9 <cjk>
	`交`: [u8(0x8C), 0xF0] // U+4EA4 <cjk>
	`佼`: [u8(0x8C), 0xF1] // U+4F7C <cjk>
	`侯`: [u8(0x8C), 0xF2] // U+4FAF <cjk>
	`候`: [u8(0x8C), 0xF3] // U+5019 <cjk>
	`倖`: [u8(0x8C), 0xF4] // U+5016 <cjk>
	`光`: [u8(0x8C), 0xF5] // U+5149 <cjk>
	`公`: [u8(0x8C), 0xF6] // U+516C <cjk>
	`功`: [u8(0x8C), 0xF7] // U+529F <cjk>
	`効`: [u8(0x8C), 0xF8] // U+52B9 <cjk>
	`勾`: [u8(0x8C), 0xF9] // U+52FE <cjk>
	`厚`: [u8(0x8C), 0xFA] // U+539A <cjk>
	`口`: [u8(0x8C), 0xFB] // U+53E3 <cjk>
	`向`: [u8(0x8C), 0xFC] // U+5411 <cjk>
	`后`: [u8(0x8D), 0x40] // U+540E <cjk>
	`喉`: [u8(0x8D), 0x41] // U+5589 <cjk>
	`坑`: [u8(0x8D), 0x42] // U+5751 <cjk>
	`垢`: [u8(0x8D), 0x43] // U+57A2 <cjk>
	`好`: [u8(0x8D), 0x44] // U+597D <cjk>
	`孔`: [u8(0x8D), 0x45] // U+5B54 <cjk>
	`孝`: [u8(0x8D), 0x46] // U+5B5D <cjk>
	`宏`: [u8(0x8D), 0x47] // U+5B8F <cjk>
	`工`: [u8(0x8D), 0x48] // U+5DE5 <cjk>
	`巧`: [u8(0x8D), 0x49] // U+5DE7 <cjk>
	`巷`: [u8(0x8D), 0x4A] // U+5DF7 <cjk>
	`幸`: [u8(0x8D), 0x4B] // U+5E78 <cjk>
	`広`: [u8(0x8D), 0x4C] // U+5E83 <cjk>
	`庚`: [u8(0x8D), 0x4D] // U+5E9A <cjk>
	`康`: [u8(0x8D), 0x4E] // U+5EB7 <cjk>
	`弘`: [u8(0x8D), 0x4F] // U+5F18 <cjk>
	`恒`: [u8(0x8D), 0x50] // U+6052 <cjk>
	`慌`: [u8(0x8D), 0x51] // U+614C <cjk>
	`抗`: [u8(0x8D), 0x52] // U+6297 <cjk>
	`拘`: [u8(0x8D), 0x53] // U+62D8 <cjk>
	`控`: [u8(0x8D), 0x54] // U+63A7 <cjk>
	`攻`: [u8(0x8D), 0x55] // U+653B <cjk>
	`昂`: [u8(0x8D), 0x56] // U+6602 <cjk>
	`晃`: [u8(0x8D), 0x57] // U+6643 <cjk>
	`更`: [u8(0x8D), 0x58] // U+66F4 <cjk>
	`杭`: [u8(0x8D), 0x59] // U+676D <cjk>
	`校`: [u8(0x8D), 0x5A] // U+6821 <cjk>
	`梗`: [u8(0x8D), 0x5B] // U+6897 <cjk>
	`構`: [u8(0x8D), 0x5C] // U+69CB <cjk>
	`江`: [u8(0x8D), 0x5D] // U+6C5F <cjk>
	`洪`: [u8(0x8D), 0x5E] // U+6D2A <cjk>
	`浩`: [u8(0x8D), 0x5F] // U+6D69 <cjk>
	`港`: [u8(0x8D), 0x60] // U+6E2F <cjk>
	`溝`: [u8(0x8D), 0x61] // U+6E9D <cjk>
	`甲`: [u8(0x8D), 0x62] // U+7532 <cjk>
	`皇`: [u8(0x8D), 0x63] // U+7687 <cjk>
	`硬`: [u8(0x8D), 0x64] // U+786C <cjk>
	`稿`: [u8(0x8D), 0x65] // U+7A3F <cjk>
	`糠`: [u8(0x8D), 0x66] // U+7CE0 <cjk>
	`紅`: [u8(0x8D), 0x67] // U+7D05 <cjk>
	`紘`: [u8(0x8D), 0x68] // U+7D18 <cjk>
	`絞`: [u8(0x8D), 0x69] // U+7D5E <cjk>
	`綱`: [u8(0x8D), 0x6A] // U+7DB1 <cjk>
	`耕`: [u8(0x8D), 0x6B] // U+8015 <cjk>
	`考`: [u8(0x8D), 0x6C] // U+8003 <cjk>
	`肯`: [u8(0x8D), 0x6D] // U+80AF <cjk>
	`肱`: [u8(0x8D), 0x6E] // U+80B1 <cjk>
	`腔`: [u8(0x8D), 0x6F] // U+8154 <cjk>
	`膏`: [u8(0x8D), 0x70] // U+818F <cjk>
	`航`: [u8(0x8D), 0x71] // U+822A <cjk>
	`荒`: [u8(0x8D), 0x72] // U+8352 <cjk>
	`行`: [u8(0x8D), 0x73] // U+884C <cjk>
	`衡`: [u8(0x8D), 0x74] // U+8861 <cjk>
	`講`: [u8(0x8D), 0x75] // U+8B1B <cjk>
	`貢`: [u8(0x8D), 0x76] // U+8CA2 <cjk>
	`購`: [u8(0x8D), 0x77] // U+8CFC <cjk>
	`郊`: [u8(0x8D), 0x78] // U+90CA <cjk>
	`酵`: [u8(0x8D), 0x79] // U+9175 <cjk>
	`鉱`: [u8(0x8D), 0x7A] // U+9271 <cjk>
	`砿`: [u8(0x8D), 0x7B] // U+783F <cjk>
	`鋼`: [u8(0x8D), 0x7C] // U+92FC <cjk>
	`閤`: [u8(0x8D), 0x7D] // U+95A4 <cjk>
	`降`: [u8(0x8D), 0x7E] // U+964D <cjk>
	`項`: [u8(0x8D), 0x80] // U+9805 <cjk>
	`香`: [u8(0x8D), 0x81] // U+9999 <cjk>
	`高`: [u8(0x8D), 0x82] // U+9AD8 <cjk>
	`鴻`: [u8(0x8D), 0x83] // U+9D3B <cjk>
	`剛`: [u8(0x8D), 0x84] // U+525B <cjk>
	`劫`: [u8(0x8D), 0x85] // U+52AB <cjk>
	`号`: [u8(0x8D), 0x86] // U+53F7 <cjk>
	`合`: [u8(0x8D), 0x87] // U+5408 <cjk>
	`壕`: [u8(0x8D), 0x88] // U+58D5 <cjk>
	`拷`: [u8(0x8D), 0x89] // U+62F7 <cjk>
	`濠`: [u8(0x8D), 0x8A] // U+6FE0 <cjk>
	`豪`: [u8(0x8D), 0x8B] // U+8C6A <cjk>
	`轟`: [u8(0x8D), 0x8C] // U+8F5F <cjk>
	`麹`: [u8(0x8D), 0x8D] // U+9EB9 <cjk>
	`克`: [u8(0x8D), 0x8E] // U+514B <cjk>
	`刻`: [u8(0x8D), 0x8F] // U+523B <cjk>
	`告`: [u8(0x8D), 0x90] // U+544A <cjk>
	`国`: [u8(0x8D), 0x91] // U+56FD <cjk>
	`穀`: [u8(0x8D), 0x92] // U+7A40 <cjk>
	`酷`: [u8(0x8D), 0x93] // U+9177 <cjk>
	`鵠`: [u8(0x8D), 0x94] // U+9D60 <cjk>
	`黒`: [u8(0x8D), 0x95] // U+9ED2 <cjk>
	`獄`: [u8(0x8D), 0x96] // U+7344 <cjk>
	`漉`: [u8(0x8D), 0x97] // U+6F09 <cjk>
	`腰`: [u8(0x8D), 0x98] // U+8170 <cjk>
	`甑`: [u8(0x8D), 0x99] // U+7511 <cjk>
	`忽`: [u8(0x8D), 0x9A] // U+5FFD <cjk>
	`惚`: [u8(0x8D), 0x9B] // U+60DA <cjk>
	`骨`: [u8(0x8D), 0x9C] // U+9AA8 <cjk>
	`狛`: [u8(0x8D), 0x9D] // U+72DB <cjk>
	`込`: [u8(0x8D), 0x9E] // U+8FBC <cjk>
	`此`: [u8(0x8D), 0x9F] // U+6B64 <cjk>
	`頃`: [u8(0x8D), 0xA0] // U+9803 <cjk>
	`今`: [u8(0x8D), 0xA1] // U+4ECA <cjk>
	`困`: [u8(0x8D), 0xA2] // U+56F0 <cjk>
	`坤`: [u8(0x8D), 0xA3] // U+5764 <cjk>
	`墾`: [u8(0x8D), 0xA4] // U+58BE <cjk>
	`婚`: [u8(0x8D), 0xA5] // U+5A5A <cjk>
	`恨`: [u8(0x8D), 0xA6] // U+6068 <cjk>
	`懇`: [u8(0x8D), 0xA7] // U+61C7 <cjk>
	`昏`: [u8(0x8D), 0xA8] // U+660F <cjk>
	`昆`: [u8(0x8D), 0xA9] // U+6606 <cjk>
	`根`: [u8(0x8D), 0xAA] // U+6839 <cjk>
	`梱`: [u8(0x8D), 0xAB] // U+68B1 <cjk>
	`混`: [u8(0x8D), 0xAC] // U+6DF7 <cjk>
	`痕`: [u8(0x8D), 0xAD] // U+75D5 <cjk>
	`紺`: [u8(0x8D), 0xAE] // U+7D3A <cjk>
	`艮`: [u8(0x8D), 0xAF] // U+826E <cjk>
	`魂`: [u8(0x8D), 0xB0] // U+9B42 <cjk>
	`些`: [u8(0x8D), 0xB1] // U+4E9B <cjk>
	`佐`: [u8(0x8D), 0xB2] // U+4F50 <cjk>
	`叉`: [u8(0x8D), 0xB3] // U+53C9 <cjk>
	`唆`: [u8(0x8D), 0xB4] // U+5506 <cjk>
	`嵯`: [u8(0x8D), 0xB5] // U+5D6F <cjk>
	`左`: [u8(0x8D), 0xB6] // U+5DE6 <cjk>
	`差`: [u8(0x8D), 0xB7] // U+5DEE <cjk>
	`査`: [u8(0x8D), 0xB8] // U+67FB <cjk>
	`沙`: [u8(0x8D), 0xB9] // U+6C99 <cjk>
	`瑳`: [u8(0x8D), 0xBA] // U+7473 <cjk>
	`砂`: [u8(0x8D), 0xBB] // U+7802 <cjk>
	`詐`: [u8(0x8D), 0xBC] // U+8A50 <cjk>
	`鎖`: [u8(0x8D), 0xBD] // U+9396 <cjk>
	`裟`: [u8(0x8D), 0xBE] // U+88DF <cjk>
	`坐`: [u8(0x8D), 0xBF] // U+5750 <cjk>
	`座`: [u8(0x8D), 0xC0] // U+5EA7 <cjk>
	`挫`: [u8(0x8D), 0xC1] // U+632B <cjk>
	`債`: [u8(0x8D), 0xC2] // U+50B5 <cjk>
	`催`: [u8(0x8D), 0xC3] // U+50AC <cjk>
	`再`: [u8(0x8D), 0xC4] // U+518D <cjk>
	`最`: [u8(0x8D), 0xC5] // U+6700 <cjk>
	`哉`: [u8(0x8D), 0xC6] // U+54C9 <cjk>
	`塞`: [u8(0x8D), 0xC7] // U+585E <cjk>
	`妻`: [u8(0x8D), 0xC8] // U+59BB <cjk>
	`宰`: [u8(0x8D), 0xC9] // U+5BB0 <cjk>
	`彩`: [u8(0x8D), 0xCA] // U+5F69 <cjk>
	`才`: [u8(0x8D), 0xCB] // U+624D <cjk>
	`採`: [u8(0x8D), 0xCC] // U+63A1 <cjk>
	`栽`: [u8(0x8D), 0xCD] // U+683D <cjk>
	`歳`: [u8(0x8D), 0xCE] // U+6B73 <cjk>
	`済`: [u8(0x8D), 0xCF] // U+6E08 <cjk>
	`災`: [u8(0x8D), 0xD0] // U+707D <cjk>
	`采`: [u8(0x8D), 0xD1] // U+91C7 <cjk>
	`犀`: [u8(0x8D), 0xD2] // U+7280 <cjk>
	`砕`: [u8(0x8D), 0xD3] // U+7815 <cjk>
	`砦`: [u8(0x8D), 0xD4] // U+7826 <cjk>
	`祭`: [u8(0x8D), 0xD5] // U+796D <cjk>
	`斎`: [u8(0x8D), 0xD6] // U+658E <cjk>
	`細`: [u8(0x8D), 0xD7] // U+7D30 <cjk>
	`菜`: [u8(0x8D), 0xD8] // U+83DC <cjk>
	`裁`: [u8(0x8D), 0xD9] // U+88C1 <cjk>
	`載`: [u8(0x8D), 0xDA] // U+8F09 <cjk>
	`際`: [u8(0x8D), 0xDB] // U+969B <cjk>
	`剤`: [u8(0x8D), 0xDC] // U+5264 <cjk>
	`在`: [u8(0x8D), 0xDD] // U+5728 <cjk>
	`材`: [u8(0x8D), 0xDE] // U+6750 <cjk>
	`罪`: [u8(0x8D), 0xDF] // U+7F6A <cjk>
	`財`: [u8(0x8D), 0xE0] // U+8CA1 <cjk>
	`冴`: [u8(0x8D), 0xE1] // U+51B4 <cjk>
	`坂`: [u8(0x8D), 0xE2] // U+5742 <cjk>
	`阪`: [u8(0x8D), 0xE3] // U+962A <cjk>
	`堺`: [u8(0x8D), 0xE4] // U+583A <cjk>
	`榊`: [u8(0x8D), 0xE5] // U+698A <cjk>
	`肴`: [u8(0x8D), 0xE6] // U+80B4 <cjk>
	`咲`: [u8(0x8D), 0xE7] // U+54B2 <cjk>
	`崎`: [u8(0x8D), 0xE8] // U+5D0E <cjk>
	`埼`: [u8(0x8D), 0xE9] // U+57FC <cjk>
	`碕`: [u8(0x8D), 0xEA] // U+7895 <cjk>
	`鷺`: [u8(0x8D), 0xEB] // U+9DFA <cjk>
	`作`: [u8(0x8D), 0xEC] // U+4F5C <cjk>
	`削`: [u8(0x8D), 0xED] // U+524A <cjk>
	`咋`: [u8(0x8D), 0xEE] // U+548B <cjk>
	`搾`: [u8(0x8D), 0xEF] // U+643E <cjk>
	`昨`: [u8(0x8D), 0xF0] // U+6628 <cjk>
	`朔`: [u8(0x8D), 0xF1] // U+6714 <cjk>
	`柵`: [u8(0x8D), 0xF2] // U+67F5 <cjk>
	`窄`: [u8(0x8D), 0xF3] // U+7A84 <cjk>
	`策`: [u8(0x8D), 0xF4] // U+7B56 <cjk>
	`索`: [u8(0x8D), 0xF5] // U+7D22 <cjk>
	`錯`: [u8(0x8D), 0xF6] // U+932F <cjk>
	`桜`: [u8(0x8D), 0xF7] // U+685C <cjk>
	`鮭`: [u8(0x8D), 0xF8] // U+9BAD <cjk>
	`笹`: [u8(0x8D), 0xF9] // U+7B39 <cjk>
	`匙`: [u8(0x8D), 0xFA] // U+5319 <cjk>
	`冊`: [u8(0x8D), 0xFB] // U+518A <cjk>
	`刷`: [u8(0x8D), 0xFC] // U+5237 <cjk>
	`察`: [u8(0x8E), 0x40] // U+5BDF <cjk>
	`拶`: [u8(0x8E), 0x41] // U+62F6 <cjk>
	`撮`: [u8(0x8E), 0x42] // U+64AE <cjk>
	`擦`: [u8(0x8E), 0x43] // U+64E6 <cjk>
	`札`: [u8(0x8E), 0x44] // U+672D <cjk>
	`殺`: [u8(0x8E), 0x45] // U+6BBA <cjk>
	`薩`: [u8(0x8E), 0x46] // U+85A9 <cjk>
	`雑`: [u8(0x8E), 0x47] // U+96D1 <cjk>
	`皐`: [u8(0x8E), 0x48] // U+7690 <cjk>
	`鯖`: [u8(0x8E), 0x49] // U+9BD6 <cjk>
	`捌`: [u8(0x8E), 0x4A] // U+634C <cjk>
	`錆`: [u8(0x8E), 0x4B] // U+9306 <cjk>
	`鮫`: [u8(0x8E), 0x4C] // U+9BAB <cjk>
	`皿`: [u8(0x8E), 0x4D] // U+76BF <cjk>
	`晒`: [u8(0x8E), 0x4E] // U+6652 <cjk>
	`三`: [u8(0x8E), 0x4F] // U+4E09 <cjk>
	`傘`: [u8(0x8E), 0x50] // U+5098 <cjk>
	`参`: [u8(0x8E), 0x51] // U+53C2 <cjk>
	`山`: [u8(0x8E), 0x52] // U+5C71 <cjk>
	`惨`: [u8(0x8E), 0x53] // U+60E8 <cjk>
	`撒`: [u8(0x8E), 0x54] // U+6492 <cjk>
	`散`: [u8(0x8E), 0x55] // U+6563 <cjk>
	`桟`: [u8(0x8E), 0x56] // U+685F <cjk>
	`燦`: [u8(0x8E), 0x57] // U+71E6 <cjk>
	`珊`: [u8(0x8E), 0x58] // U+73CA <cjk>
	`産`: [u8(0x8E), 0x59] // U+7523 <cjk>
	`算`: [u8(0x8E), 0x5A] // U+7B97 <cjk>
	`纂`: [u8(0x8E), 0x5B] // U+7E82 <cjk>
	`蚕`: [u8(0x8E), 0x5C] // U+8695 <cjk>
	`讃`: [u8(0x8E), 0x5D] // U+8B83 <cjk>
	`賛`: [u8(0x8E), 0x5E] // U+8CDB <cjk>
	`酸`: [u8(0x8E), 0x5F] // U+9178 <cjk>
	`餐`: [u8(0x8E), 0x60] // U+9910 <cjk>
	`斬`: [u8(0x8E), 0x61] // U+65AC <cjk>
	`暫`: [u8(0x8E), 0x62] // U+66AB <cjk>
	`残`: [u8(0x8E), 0x63] // U+6B8B <cjk>
	`仕`: [u8(0x8E), 0x64] // U+4ED5 <cjk>
	`仔`: [u8(0x8E), 0x65] // U+4ED4 <cjk>
	`伺`: [u8(0x8E), 0x66] // U+4F3A <cjk>
	`使`: [u8(0x8E), 0x67] // U+4F7F <cjk>
	`刺`: [u8(0x8E), 0x68] // U+523A <cjk>
	`司`: [u8(0x8E), 0x69] // U+53F8 <cjk>
	`史`: [u8(0x8E), 0x6A] // U+53F2 <cjk>
	`嗣`: [u8(0x8E), 0x6B] // U+55E3 <cjk>
	`四`: [u8(0x8E), 0x6C] // U+56DB <cjk>
	`士`: [u8(0x8E), 0x6D] // U+58EB <cjk>
	`始`: [u8(0x8E), 0x6E] // U+59CB <cjk>
	`姉`: [u8(0x8E), 0x6F] // U+59C9 <cjk>
	`姿`: [u8(0x8E), 0x70] // U+59FF <cjk>
	`子`: [u8(0x8E), 0x71] // U+5B50 <cjk>
	`屍`: [u8(0x8E), 0x72] // U+5C4D <cjk>
	`市`: [u8(0x8E), 0x73] // U+5E02 <cjk>
	`師`: [u8(0x8E), 0x74] // U+5E2B <cjk>
	`志`: [u8(0x8E), 0x75] // U+5FD7 <cjk>
	`思`: [u8(0x8E), 0x76] // U+601D <cjk>
	`指`: [u8(0x8E), 0x77] // U+6307 <cjk>
	`支`: [u8(0x8E), 0x78] // U+652F <cjk>
	`孜`: [u8(0x8E), 0x79] // U+5B5C <cjk>
	`斯`: [u8(0x8E), 0x7A] // U+65AF <cjk>
	`施`: [u8(0x8E), 0x7B] // U+65BD <cjk>
	`旨`: [u8(0x8E), 0x7C] // U+65E8 <cjk>
	`枝`: [u8(0x8E), 0x7D] // U+679D <cjk>
	`止`: [u8(0x8E), 0x7E] // U+6B62 <cjk>
	`死`: [u8(0x8E), 0x80] // U+6B7B <cjk>
	`氏`: [u8(0x8E), 0x81] // U+6C0F <cjk>
	`獅`: [u8(0x8E), 0x82] // U+7345 <cjk>
	`祉`: [u8(0x8E), 0x83] // U+7949 <cjk>
	`私`: [u8(0x8E), 0x84] // U+79C1 <cjk>
	`糸`: [u8(0x8E), 0x85] // U+7CF8 <cjk>
	`紙`: [u8(0x8E), 0x86] // U+7D19 <cjk>
	`紫`: [u8(0x8E), 0x87] // U+7D2B <cjk>
	`肢`: [u8(0x8E), 0x88] // U+80A2 <cjk>
	`脂`: [u8(0x8E), 0x89] // U+8102 <cjk>
	`至`: [u8(0x8E), 0x8A] // U+81F3 <cjk>
	`視`: [u8(0x8E), 0x8B] // U+8996 <cjk>
	`詞`: [u8(0x8E), 0x8C] // U+8A5E <cjk>
	`詩`: [u8(0x8E), 0x8D] // U+8A69 <cjk>
	`試`: [u8(0x8E), 0x8E] // U+8A66 <cjk>
	`誌`: [u8(0x8E), 0x8F] // U+8A8C <cjk>
	`諮`: [u8(0x8E), 0x90] // U+8AEE <cjk>
	`資`: [u8(0x8E), 0x91] // U+8CC7 <cjk>
	`賜`: [u8(0x8E), 0x92] // U+8CDC <cjk>
	`雌`: [u8(0x8E), 0x93] // U+96CC <cjk>
	`飼`: [u8(0x8E), 0x94] // U+98FC <cjk>
	`歯`: [u8(0x8E), 0x95] // U+6B6F <cjk>
	`事`: [u8(0x8E), 0x96] // U+4E8B <cjk>
	`似`: [u8(0x8E), 0x97] // U+4F3C <cjk>
	`侍`: [u8(0x8E), 0x98] // U+4F8D <cjk>
	`児`: [u8(0x8E), 0x99] // U+5150 <cjk>
	`字`: [u8(0x8E), 0x9A] // U+5B57 <cjk>
	`寺`: [u8(0x8E), 0x9B] // U+5BFA <cjk>
	`慈`: [u8(0x8E), 0x9C] // U+6148 <cjk>
	`持`: [u8(0x8E), 0x9D] // U+6301 <cjk>
	`時`: [u8(0x8E), 0x9E] // U+6642 <cjk>
	`次`: [u8(0x8E), 0x9F] // U+6B21 <cjk>
	`滋`: [u8(0x8E), 0xA0] // U+6ECB <cjk>
	`治`: [u8(0x8E), 0xA1] // U+6CBB <cjk>
	`爾`: [u8(0x8E), 0xA2] // U+723E <cjk>
	`璽`: [u8(0x8E), 0xA3] // U+74BD <cjk>
	`痔`: [u8(0x8E), 0xA4] // U+75D4 <cjk>
	`磁`: [u8(0x8E), 0xA5] // U+78C1 <cjk>
	`示`: [u8(0x8E), 0xA6] // U+793A <cjk>
	`而`: [u8(0x8E), 0xA7] // U+800C <cjk>
	`耳`: [u8(0x8E), 0xA8] // U+8033 <cjk>
	`自`: [u8(0x8E), 0xA9] // U+81EA <cjk>
	`蒔`: [u8(0x8E), 0xAA] // U+8494 <cjk>
	`辞`: [u8(0x8E), 0xAB] // U+8F9E <cjk>
	`汐`: [u8(0x8E), 0xAC] // U+6C50 <cjk>
	`鹿`: [u8(0x8E), 0xAD] // U+9E7F <cjk>
	`式`: [u8(0x8E), 0xAE] // U+5F0F <cjk>
	`識`: [u8(0x8E), 0xAF] // U+8B58 <cjk>
	`鴫`: [u8(0x8E), 0xB0] // U+9D2B <cjk>
	`竺`: [u8(0x8E), 0xB1] // U+7AFA <cjk>
	`軸`: [u8(0x8E), 0xB2] // U+8EF8 <cjk>
	`宍`: [u8(0x8E), 0xB3] // U+5B8D <cjk>
	`雫`: [u8(0x8E), 0xB4] // U+96EB <cjk>
	`七`: [u8(0x8E), 0xB5] // U+4E03 <cjk>
	`叱`: [u8(0x8E), 0xB6] // U+53F1 <cjk>
	`執`: [u8(0x8E), 0xB7] // U+57F7 <cjk>
	`失`: [u8(0x8E), 0xB8] // U+5931 <cjk>
	`嫉`: [u8(0x8E), 0xB9] // U+5AC9 <cjk>
	`室`: [u8(0x8E), 0xBA] // U+5BA4 <cjk>
	`悉`: [u8(0x8E), 0xBB] // U+6089 <cjk>
	`湿`: [u8(0x8E), 0xBC] // U+6E7F <cjk>
	`漆`: [u8(0x8E), 0xBD] // U+6F06 <cjk>
	`疾`: [u8(0x8E), 0xBE] // U+75BE <cjk>
	`質`: [u8(0x8E), 0xBF] // U+8CEA <cjk>
	`実`: [u8(0x8E), 0xC0] // U+5B9F <cjk>
	`蔀`: [u8(0x8E), 0xC1] // U+8500 <cjk>
	`篠`: [u8(0x8E), 0xC2] // U+7BE0 <cjk>
	`偲`: [u8(0x8E), 0xC3] // U+5072 <cjk>
	`柴`: [u8(0x8E), 0xC4] // U+67F4 <cjk>
	`芝`: [u8(0x8E), 0xC5] // U+829D <cjk>
	`屡`: [u8(0x8E), 0xC6] // U+5C61 <cjk>
	`蕊`: [u8(0x8E), 0xC7] // U+854A <cjk>
	`縞`: [u8(0x8E), 0xC8] // U+7E1E <cjk>
	`舎`: [u8(0x8E), 0xC9] // U+820E <cjk>
	`写`: [u8(0x8E), 0xCA] // U+5199 <cjk>
	`射`: [u8(0x8E), 0xCB] // U+5C04 <cjk>
	`捨`: [u8(0x8E), 0xCC] // U+6368 <cjk>
	`赦`: [u8(0x8E), 0xCD] // U+8D66 <cjk>
	`斜`: [u8(0x8E), 0xCE] // U+659C <cjk>
	`煮`: [u8(0x8E), 0xCF] // U+716E <cjk>
	`社`: [u8(0x8E), 0xD0] // U+793E <cjk>
	`紗`: [u8(0x8E), 0xD1] // U+7D17 <cjk>
	`者`: [u8(0x8E), 0xD2] // U+8005 <cjk>
	`謝`: [u8(0x8E), 0xD3] // U+8B1D <cjk>
	`車`: [u8(0x8E), 0xD4] // U+8ECA <cjk>
	`遮`: [u8(0x8E), 0xD5] // U+906E <cjk>
	`蛇`: [u8(0x8E), 0xD6] // U+86C7 <cjk>
	`邪`: [u8(0x8E), 0xD7] // U+90AA <cjk>
	`借`: [u8(0x8E), 0xD8] // U+501F <cjk>
	`勺`: [u8(0x8E), 0xD9] // U+52FA <cjk>
	`尺`: [u8(0x8E), 0xDA] // U+5C3A <cjk>
	`杓`: [u8(0x8E), 0xDB] // U+6753 <cjk>
	`灼`: [u8(0x8E), 0xDC] // U+707C <cjk>
	`爵`: [u8(0x8E), 0xDD] // U+7235 <cjk>
	`酌`: [u8(0x8E), 0xDE] // U+914C <cjk>
	`釈`: [u8(0x8E), 0xDF] // U+91C8 <cjk>
	`錫`: [u8(0x8E), 0xE0] // U+932B <cjk>
	`若`: [u8(0x8E), 0xE1] // U+82E5 <cjk>
	`寂`: [u8(0x8E), 0xE2] // U+5BC2 <cjk>
	`弱`: [u8(0x8E), 0xE3] // U+5F31 <cjk>
	`惹`: [u8(0x8E), 0xE4] // U+60F9 <cjk>
	`主`: [u8(0x8E), 0xE5] // U+4E3B <cjk>
	`取`: [u8(0x8E), 0xE6] // U+53D6 <cjk>
	`守`: [u8(0x8E), 0xE7] // U+5B88 <cjk>
	`手`: [u8(0x8E), 0xE8] // U+624B <cjk>
	`朱`: [u8(0x8E), 0xE9] // U+6731 <cjk>
	`殊`: [u8(0x8E), 0xEA] // U+6B8A <cjk>
	`狩`: [u8(0x8E), 0xEB] // U+72E9 <cjk>
	`珠`: [u8(0x8E), 0xEC] // U+73E0 <cjk>
	`種`: [u8(0x8E), 0xED] // U+7A2E <cjk>
	`腫`: [u8(0x8E), 0xEE] // U+816B <cjk>
	`趣`: [u8(0x8E), 0xEF] // U+8DA3 <cjk>
	`酒`: [u8(0x8E), 0xF0] // U+9152 <cjk>
	`首`: [u8(0x8E), 0xF1] // U+9996 <cjk>
	`儒`: [u8(0x8E), 0xF2] // U+5112 <cjk>
	`受`: [u8(0x8E), 0xF3] // U+53D7 <cjk>
	`呪`: [u8(0x8E), 0xF4] // U+546A <cjk>
	`寿`: [u8(0x8E), 0xF5] // U+5BFF <cjk>
	`授`: [u8(0x8E), 0xF6] // U+6388 <cjk>
	`樹`: [u8(0x8E), 0xF7] // U+6A39 <cjk>
	`綬`: [u8(0x8E), 0xF8] // U+7DAC <cjk>
	`需`: [u8(0x8E), 0xF9] // U+9700 <cjk>
	`囚`: [u8(0x8E), 0xFA] // U+56DA <cjk>
	`収`: [u8(0x8E), 0xFB] // U+53CE <cjk>
	`周`: [u8(0x8E), 0xFC] // U+5468 <cjk>
	`宗`: [u8(0x8F), 0x40] // U+5B97 <cjk>
	`就`: [u8(0x8F), 0x41] // U+5C31 <cjk>
	`州`: [u8(0x8F), 0x42] // U+5DDE <cjk>
	`修`: [u8(0x8F), 0x43] // U+4FEE <cjk>
	`愁`: [u8(0x8F), 0x44] // U+6101 <cjk>
	`拾`: [u8(0x8F), 0x45] // U+62FE <cjk>
	`洲`: [u8(0x8F), 0x46] // U+6D32 <cjk>
	`秀`: [u8(0x8F), 0x47] // U+79C0 <cjk>
	`秋`: [u8(0x8F), 0x48] // U+79CB <cjk>
	`終`: [u8(0x8F), 0x49] // U+7D42 <cjk>
	`繍`: [u8(0x8F), 0x4A] // U+7E4D <cjk>
	`習`: [u8(0x8F), 0x4B] // U+7FD2 <cjk>
	`臭`: [u8(0x8F), 0x4C] // U+81ED <cjk>
	`舟`: [u8(0x8F), 0x4D] // U+821F <cjk>
	`蒐`: [u8(0x8F), 0x4E] // U+8490 <cjk>
	`衆`: [u8(0x8F), 0x4F] // U+8846 <cjk>
	`襲`: [u8(0x8F), 0x50] // U+8972 <cjk>
	`讐`: [u8(0x8F), 0x51] // U+8B90 <cjk>
	`蹴`: [u8(0x8F), 0x52] // U+8E74 <cjk>
	`輯`: [u8(0x8F), 0x53] // U+8F2F <cjk>
	`週`: [u8(0x8F), 0x54] // U+9031 <cjk>
	`酋`: [u8(0x8F), 0x55] // U+914B <cjk>
	`酬`: [u8(0x8F), 0x56] // U+916C <cjk>
	`集`: [u8(0x8F), 0x57] // U+96C6 <cjk>
	`醜`: [u8(0x8F), 0x58] // U+919C <cjk>
	`什`: [u8(0x8F), 0x59] // U+4EC0 <cjk>
	`住`: [u8(0x8F), 0x5A] // U+4F4F <cjk>
	`充`: [u8(0x8F), 0x5B] // U+5145 <cjk>
	`十`: [u8(0x8F), 0x5C] // U+5341 <cjk>
	`従`: [u8(0x8F), 0x5D] // U+5F93 <cjk>
	`戎`: [u8(0x8F), 0x5E] // U+620E <cjk>
	`柔`: [u8(0x8F), 0x5F] // U+67D4 <cjk>
	`汁`: [u8(0x8F), 0x60] // U+6C41 <cjk>
	`渋`: [u8(0x8F), 0x61] // U+6E0B <cjk>
	`獣`: [u8(0x8F), 0x62] // U+7363 <cjk>
	`縦`: [u8(0x8F), 0x63] // U+7E26 <cjk>
	`重`: [u8(0x8F), 0x64] // U+91CD <cjk>
	`銃`: [u8(0x8F), 0x65] // U+9283 <cjk>
	`叔`: [u8(0x8F), 0x66] // U+53D4 <cjk>
	`夙`: [u8(0x8F), 0x67] // U+5919 <cjk>
	`宿`: [u8(0x8F), 0x68] // U+5BBF <cjk>
	`淑`: [u8(0x8F), 0x69] // U+6DD1 <cjk>
	`祝`: [u8(0x8F), 0x6A] // U+795D <cjk>
	`縮`: [u8(0x8F), 0x6B] // U+7E2E <cjk>
	`粛`: [u8(0x8F), 0x6C] // U+7C9B <cjk>
	`塾`: [u8(0x8F), 0x6D] // U+587E <cjk>
	`熟`: [u8(0x8F), 0x6E] // U+719F <cjk>
	`出`: [u8(0x8F), 0x6F] // U+51FA <cjk>
	`術`: [u8(0x8F), 0x70] // U+8853 <cjk>
	`述`: [u8(0x8F), 0x71] // U+8FF0 <cjk>
	`俊`: [u8(0x8F), 0x72] // U+4FCA <cjk>
	`峻`: [u8(0x8F), 0x73] // U+5CFB <cjk>
	`春`: [u8(0x8F), 0x74] // U+6625 <cjk>
	`瞬`: [u8(0x8F), 0x75] // U+77AC <cjk>
	`竣`: [u8(0x8F), 0x76] // U+7AE3 <cjk>
	`舜`: [u8(0x8F), 0x77] // U+821C <cjk>
	`駿`: [u8(0x8F), 0x78] // U+99FF <cjk>
	`准`: [u8(0x8F), 0x79] // U+51C6 <cjk>
	`循`: [u8(0x8F), 0x7A] // U+5FAA <cjk>
	`旬`: [u8(0x8F), 0x7B] // U+65EC <cjk>
	`楯`: [u8(0x8F), 0x7C] // U+696F <cjk>
	`殉`: [u8(0x8F), 0x7D] // U+6B89 <cjk>
	`淳`: [u8(0x8F), 0x7E] // U+6DF3 <cjk>
	`準`: [u8(0x8F), 0x80] // U+6E96 <cjk>
	`潤`: [u8(0x8F), 0x81] // U+6F64 <cjk>
	`盾`: [u8(0x8F), 0x82] // U+76FE <cjk>
	`純`: [u8(0x8F), 0x83] // U+7D14 <cjk>
	`巡`: [u8(0x8F), 0x84] // U+5DE1 <cjk>
	`遵`: [u8(0x8F), 0x85] // U+9075 <cjk>
	`醇`: [u8(0x8F), 0x86] // U+9187 <cjk>
	`順`: [u8(0x8F), 0x87] // U+9806 <cjk>
	`処`: [u8(0x8F), 0x88] // U+51E6 <cjk>
	`初`: [u8(0x8F), 0x89] // U+521D <cjk>
	`所`: [u8(0x8F), 0x8A] // U+6240 <cjk>
	`暑`: [u8(0x8F), 0x8B] // U+6691 <cjk>
	`曙`: [u8(0x8F), 0x8C] // U+66D9 <cjk>
	`渚`: [u8(0x8F), 0x8D] // U+6E1A <cjk>
	`庶`: [u8(0x8F), 0x8E] // U+5EB6 <cjk>
	`緒`: [u8(0x8F), 0x8F] // U+7DD2 <cjk>
	`署`: [u8(0x8F), 0x90] // U+7F72 <cjk>
	`書`: [u8(0x8F), 0x91] // U+66F8 <cjk>
	`薯`: [u8(0x8F), 0x92] // U+85AF <cjk>
	`藷`: [u8(0x8F), 0x93] // U+85F7 <cjk>
	`諸`: [u8(0x8F), 0x94] // U+8AF8 <cjk>
	`助`: [u8(0x8F), 0x95] // U+52A9 <cjk>
	`叙`: [u8(0x8F), 0x96] // U+53D9 <cjk>
	`女`: [u8(0x8F), 0x97] // U+5973 <cjk>
	`序`: [u8(0x8F), 0x98] // U+5E8F <cjk>
	`徐`: [u8(0x8F), 0x99] // U+5F90 <cjk>
	`恕`: [u8(0x8F), 0x9A] // U+6055 <cjk>
	`鋤`: [u8(0x8F), 0x9B] // U+92E4 <cjk>
	`除`: [u8(0x8F), 0x9C] // U+9664 <cjk>
	`傷`: [u8(0x8F), 0x9D] // U+50B7 <cjk>
	`償`: [u8(0x8F), 0x9E] // U+511F <cjk>
	`勝`: [u8(0x8F), 0x9F] // U+52DD <cjk>
	`匠`: [u8(0x8F), 0xA0] // U+5320 <cjk>
	`升`: [u8(0x8F), 0xA1] // U+5347 <cjk>
	`召`: [u8(0x8F), 0xA2] // U+53EC <cjk>
	`哨`: [u8(0x8F), 0xA3] // U+54E8 <cjk>
	`商`: [u8(0x8F), 0xA4] // U+5546 <cjk>
	`唱`: [u8(0x8F), 0xA5] // U+5531 <cjk>
	`嘗`: [u8(0x8F), 0xA6] // U+5617 <cjk>
	`奨`: [u8(0x8F), 0xA7] // U+5968 <cjk>
	`妾`: [u8(0x8F), 0xA8] // U+59BE <cjk>
	`娼`: [u8(0x8F), 0xA9] // U+5A3C <cjk>
	`宵`: [u8(0x8F), 0xAA] // U+5BB5 <cjk>
	`将`: [u8(0x8F), 0xAB] // U+5C06 <cjk>
	`小`: [u8(0x8F), 0xAC] // U+5C0F <cjk>
	`少`: [u8(0x8F), 0xAD] // U+5C11 <cjk>
	`尚`: [u8(0x8F), 0xAE] // U+5C1A <cjk>
	`庄`: [u8(0x8F), 0xAF] // U+5E84 <cjk>
	`床`: [u8(0x8F), 0xB0] // U+5E8A <cjk>
	`廠`: [u8(0x8F), 0xB1] // U+5EE0 <cjk>
	`彰`: [u8(0x8F), 0xB2] // U+5F70 <cjk>
	`承`: [u8(0x8F), 0xB3] // U+627F <cjk>
	`抄`: [u8(0x8F), 0xB4] // U+6284 <cjk>
	`招`: [u8(0x8F), 0xB5] // U+62DB <cjk>
	`掌`: [u8(0x8F), 0xB6] // U+638C <cjk>
	`捷`: [u8(0x8F), 0xB7] // U+6377 <cjk>
	`昇`: [u8(0x8F), 0xB8] // U+6607 <cjk>
	`昌`: [u8(0x8F), 0xB9] // U+660C <cjk>
	`昭`: [u8(0x8F), 0xBA] // U+662D <cjk>
	`晶`: [u8(0x8F), 0xBB] // U+6676 <cjk>
	`松`: [u8(0x8F), 0xBC] // U+677E <cjk>
	`梢`: [u8(0x8F), 0xBD] // U+68A2 <cjk>
	`樟`: [u8(0x8F), 0xBE] // U+6A1F <cjk>
	`樵`: [u8(0x8F), 0xBF] // U+6A35 <cjk>
	`沼`: [u8(0x8F), 0xC0] // U+6CBC <cjk>
	`消`: [u8(0x8F), 0xC1] // U+6D88 <cjk>
	`渉`: [u8(0x8F), 0xC2] // U+6E09 <cjk>
	`湘`: [u8(0x8F), 0xC3] // U+6E58 <cjk>
	`焼`: [u8(0x8F), 0xC4] // U+713C <cjk>
	`焦`: [u8(0x8F), 0xC5] // U+7126 <cjk>
	`照`: [u8(0x8F), 0xC6] // U+7167 <cjk>
	`症`: [u8(0x8F), 0xC7] // U+75C7 <cjk>
	`省`: [u8(0x8F), 0xC8] // U+7701 <cjk>
	`硝`: [u8(0x8F), 0xC9] // U+785D <cjk>
	`礁`: [u8(0x8F), 0xCA] // U+7901 <cjk>
	`祥`: [u8(0x8F), 0xCB] // U+7965 <cjk>
	`称`: [u8(0x8F), 0xCC] // U+79F0 <cjk>
	`章`: [u8(0x8F), 0xCD] // U+7AE0 <cjk>
	`笑`: [u8(0x8F), 0xCE] // U+7B11 <cjk>
	`粧`: [u8(0x8F), 0xCF] // U+7CA7 <cjk>
	`紹`: [u8(0x8F), 0xD0] // U+7D39 <cjk>
	`肖`: [u8(0x8F), 0xD1] // U+8096 <cjk>
	`菖`: [u8(0x8F), 0xD2] // U+83D6 <cjk>
	`蒋`: [u8(0x8F), 0xD3] // U+848B <cjk>
	`蕉`: [u8(0x8F), 0xD4] // U+8549 <cjk>
	`衝`: [u8(0x8F), 0xD5] // U+885D <cjk>
	`裳`: [u8(0x8F), 0xD6] // U+88F3 <cjk>
	`訟`: [u8(0x8F), 0xD7] // U+8A1F <cjk>
	`証`: [u8(0x8F), 0xD8] // U+8A3C <cjk>
	`詔`: [u8(0x8F), 0xD9] // U+8A54 <cjk>
	`詳`: [u8(0x8F), 0xDA] // U+8A73 <cjk>
	`象`: [u8(0x8F), 0xDB] // U+8C61 <cjk>
	`賞`: [u8(0x8F), 0xDC] // U+8CDE <cjk>
	`醤`: [u8(0x8F), 0xDD] // U+91A4 <cjk>
	`鉦`: [u8(0x8F), 0xDE] // U+9266 <cjk>
	`鍾`: [u8(0x8F), 0xDF] // U+937E <cjk>
	`鐘`: [u8(0x8F), 0xE0] // U+9418 <cjk>
	`障`: [u8(0x8F), 0xE1] // U+969C <cjk>
	`鞘`: [u8(0x8F), 0xE2] // U+9798 <cjk>
	`上`: [u8(0x8F), 0xE3] // U+4E0A <cjk>
	`丈`: [u8(0x8F), 0xE4] // U+4E08 <cjk>
	`丞`: [u8(0x8F), 0xE5] // U+4E1E <cjk>
	`乗`: [u8(0x8F), 0xE6] // U+4E57 <cjk>
	`冗`: [u8(0x8F), 0xE7] // U+5197 <cjk>
	`剰`: [u8(0x8F), 0xE8] // U+5270 <cjk>
	`城`: [u8(0x8F), 0xE9] // U+57CE <cjk>
	`場`: [u8(0x8F), 0xEA] // U+5834 <cjk>
	`壌`: [u8(0x8F), 0xEB] // U+58CC <cjk>
	`嬢`: [u8(0x8F), 0xEC] // U+5B22 <cjk>
	`常`: [u8(0x8F), 0xED] // U+5E38 <cjk>
	`情`: [u8(0x8F), 0xEE] // U+60C5 <cjk>
	`擾`: [u8(0x8F), 0xEF] // U+64FE <cjk>
	`条`: [u8(0x8F), 0xF0] // U+6761 <cjk>
	`杖`: [u8(0x8F), 0xF1] // U+6756 <cjk>
	`浄`: [u8(0x8F), 0xF2] // U+6D44 <cjk>
	`状`: [u8(0x8F), 0xF3] // U+72B6 <cjk>
	`畳`: [u8(0x8F), 0xF4] // U+7573 <cjk>
	`穣`: [u8(0x8F), 0xF5] // U+7A63 <cjk>
	`蒸`: [u8(0x8F), 0xF6] // U+84B8 <cjk>
	`譲`: [u8(0x8F), 0xF7] // U+8B72 <cjk>
	`醸`: [u8(0x8F), 0xF8] // U+91B8 <cjk>
	`錠`: [u8(0x8F), 0xF9] // U+9320 <cjk>
	`嘱`: [u8(0x8F), 0xFA] // U+5631 <cjk>
	`埴`: [u8(0x8F), 0xFB] // U+57F4 <cjk>
	`飾`: [u8(0x8F), 0xFC] // U+98FE <cjk>
	`拭`: [u8(0x90), 0x40] // U+62ED <cjk>
	`植`: [u8(0x90), 0x41] // U+690D <cjk>
	`殖`: [u8(0x90), 0x42] // U+6B96 <cjk>
	`燭`: [u8(0x90), 0x43] // U+71ED <cjk>
	`織`: [u8(0x90), 0x44] // U+7E54 <cjk>
	`職`: [u8(0x90), 0x45] // U+8077 <cjk>
	`色`: [u8(0x90), 0x46] // U+8272 <cjk>
	`触`: [u8(0x90), 0x47] // U+89E6 <cjk>
	`食`: [u8(0x90), 0x48] // U+98DF <cjk>
	`蝕`: [u8(0x90), 0x49] // U+8755 <cjk>
	`辱`: [u8(0x90), 0x4A] // U+8FB1 <cjk>
	`尻`: [u8(0x90), 0x4B] // U+5C3B <cjk>
	`伸`: [u8(0x90), 0x4C] // U+4F38 <cjk>
	`信`: [u8(0x90), 0x4D] // U+4FE1 <cjk>
	`侵`: [u8(0x90), 0x4E] // U+4FB5 <cjk>
	`唇`: [u8(0x90), 0x4F] // U+5507 <cjk>
	`娠`: [u8(0x90), 0x50] // U+5A20 <cjk>
	`寝`: [u8(0x90), 0x51] // U+5BDD <cjk>
	`審`: [u8(0x90), 0x52] // U+5BE9 <cjk>
	`心`: [u8(0x90), 0x53] // U+5FC3 <cjk>
	`慎`: [u8(0x90), 0x54] // U+614E <cjk>
	`振`: [u8(0x90), 0x55] // U+632F <cjk>
	`新`: [u8(0x90), 0x56] // U+65B0 <cjk>
	`晋`: [u8(0x90), 0x57] // U+664B <cjk>
	`森`: [u8(0x90), 0x58] // U+68EE <cjk>
	`榛`: [u8(0x90), 0x59] // U+699B <cjk>
	`浸`: [u8(0x90), 0x5A] // U+6D78 <cjk>
	`深`: [u8(0x90), 0x5B] // U+6DF1 <cjk>
	`申`: [u8(0x90), 0x5C] // U+7533 <cjk>
	`疹`: [u8(0x90), 0x5D] // U+75B9 <cjk>
	`真`: [u8(0x90), 0x5E] // U+771F <cjk>
	`神`: [u8(0x90), 0x5F] // U+795E <cjk>
	`秦`: [u8(0x90), 0x60] // U+79E6 <cjk>
	`紳`: [u8(0x90), 0x61] // U+7D33 <cjk>
	`臣`: [u8(0x90), 0x62] // U+81E3 <cjk>
	`芯`: [u8(0x90), 0x63] // U+82AF <cjk>
	`薪`: [u8(0x90), 0x64] // U+85AA <cjk>
	`親`: [u8(0x90), 0x65] // U+89AA <cjk>
	`診`: [u8(0x90), 0x66] // U+8A3A <cjk>
	`身`: [u8(0x90), 0x67] // U+8EAB <cjk>
	`辛`: [u8(0x90), 0x68] // U+8F9B <cjk>
	`進`: [u8(0x90), 0x69] // U+9032 <cjk>
	`針`: [u8(0x90), 0x6A] // U+91DD <cjk>
	`震`: [u8(0x90), 0x6B] // U+9707 <cjk>
	`人`: [u8(0x90), 0x6C] // U+4EBA <cjk>
	`仁`: [u8(0x90), 0x6D] // U+4EC1 <cjk>
	`刃`: [u8(0x90), 0x6E] // U+5203 <cjk>
	`塵`: [u8(0x90), 0x6F] // U+5875 <cjk>
	`壬`: [u8(0x90), 0x70] // U+58EC <cjk>
	`尋`: [u8(0x90), 0x71] // U+5C0B <cjk>
	`甚`: [u8(0x90), 0x72] // U+751A <cjk>
	`尽`: [u8(0x90), 0x73] // U+5C3D <cjk>
	`腎`: [u8(0x90), 0x74] // U+814E <cjk>
	`訊`: [u8(0x90), 0x75] // U+8A0A <cjk>
	`迅`: [u8(0x90), 0x76] // U+8FC5 <cjk>
	`陣`: [u8(0x90), 0x77] // U+9663 <cjk>
	`靭`: [u8(0x90), 0x78] // U+976D <cjk>
	`笥`: [u8(0x90), 0x79] // U+7B25 <cjk>
	`諏`: [u8(0x90), 0x7A] // U+8ACF <cjk>
	`須`: [u8(0x90), 0x7B] // U+9808 <cjk>
	`酢`: [u8(0x90), 0x7C] // U+9162 <cjk>
	`図`: [u8(0x90), 0x7D] // U+56F3 <cjk>
	`厨`: [u8(0x90), 0x7E] // U+53A8 <cjk>
	`逗`: [u8(0x90), 0x80] // U+9017 <cjk>
	`吹`: [u8(0x90), 0x81] // U+5439 <cjk>
	`垂`: [u8(0x90), 0x82] // U+5782 <cjk>
	`帥`: [u8(0x90), 0x83] // U+5E25 <cjk>
	`推`: [u8(0x90), 0x84] // U+63A8 <cjk>
	`水`: [u8(0x90), 0x85] // U+6C34 <cjk>
	`炊`: [u8(0x90), 0x86] // U+708A <cjk>
	`睡`: [u8(0x90), 0x87] // U+7761 <cjk>
	`粋`: [u8(0x90), 0x88] // U+7C8B <cjk>
	`翠`: [u8(0x90), 0x89] // U+7FE0 <cjk>
	`衰`: [u8(0x90), 0x8A] // U+8870 <cjk>
	`遂`: [u8(0x90), 0x8B] // U+9042 <cjk>
	`酔`: [u8(0x90), 0x8C] // U+9154 <cjk>
	`錐`: [u8(0x90), 0x8D] // U+9310 <cjk>
	`錘`: [u8(0x90), 0x8E] // U+9318 <cjk>
	`随`: [u8(0x90), 0x8F] // U+968F <cjk>
	`瑞`: [u8(0x90), 0x90] // U+745E <cjk>
	`髄`: [u8(0x90), 0x91] // U+9AC4 <cjk>
	`崇`: [u8(0x90), 0x92] // U+5D07 <cjk>
	`嵩`: [u8(0x90), 0x93] // U+5D69 <cjk>
	`数`: [u8(0x90), 0x94] // U+6570 <cjk>
	`枢`: [u8(0x90), 0x95] // U+67A2 <cjk>
	`趨`: [u8(0x90), 0x96] // U+8DA8 <cjk>
	`雛`: [u8(0x90), 0x97] // U+96DB <cjk>
	`据`: [u8(0x90), 0x98] // U+636E <cjk>
	`杉`: [u8(0x90), 0x99] // U+6749 <cjk>
	`椙`: [u8(0x90), 0x9A] // U+6919 <cjk>
	`菅`: [u8(0x90), 0x9B] // U+83C5 <cjk>
	`頗`: [u8(0x90), 0x9C] // U+9817 <cjk>
	`雀`: [u8(0x90), 0x9D] // U+96C0 <cjk>
	`裾`: [u8(0x90), 0x9E] // U+88FE <cjk>
	`澄`: [u8(0x90), 0x9F] // U+6F84 <cjk>
	`摺`: [u8(0x90), 0xA0] // U+647A <cjk>
	`寸`: [u8(0x90), 0xA1] // U+5BF8 <cjk>
	`世`: [u8(0x90), 0xA2] // U+4E16 <cjk>
	`瀬`: [u8(0x90), 0xA3] // U+702C <cjk>
	`畝`: [u8(0x90), 0xA4] // U+755D <cjk>
	`是`: [u8(0x90), 0xA5] // U+662F <cjk>
	`凄`: [u8(0x90), 0xA6] // U+51C4 <cjk>
	`制`: [u8(0x90), 0xA7] // U+5236 <cjk>
	`勢`: [u8(0x90), 0xA8] // U+52E2 <cjk>
	`姓`: [u8(0x90), 0xA9] // U+59D3 <cjk>
	`征`: [u8(0x90), 0xAA] // U+5F81 <cjk>
	`性`: [u8(0x90), 0xAB] // U+6027 <cjk>
	`成`: [u8(0x90), 0xAC] // U+6210 <cjk>
	`政`: [u8(0x90), 0xAD] // U+653F <cjk>
	`整`: [u8(0x90), 0xAE] // U+6574 <cjk>
	`星`: [u8(0x90), 0xAF] // U+661F <cjk>
	`晴`: [u8(0x90), 0xB0] // U+6674 <cjk>
	`棲`: [u8(0x90), 0xB1] // U+68F2 <cjk>
	`栖`: [u8(0x90), 0xB2] // U+6816 <cjk>
	`正`: [u8(0x90), 0xB3] // U+6B63 <cjk>
	`清`: [u8(0x90), 0xB4] // U+6E05 <cjk>
	`牲`: [u8(0x90), 0xB5] // U+7272 <cjk>
	`生`: [u8(0x90), 0xB6] // U+751F <cjk>
	`盛`: [u8(0x90), 0xB7] // U+76DB <cjk>
	`精`: [u8(0x90), 0xB8] // U+7CBE <cjk>
	`聖`: [u8(0x90), 0xB9] // U+8056 <cjk>
	`声`: [u8(0x90), 0xBA] // U+58F0 <cjk>
	`製`: [u8(0x90), 0xBB] // U+88FD <cjk>
	`西`: [u8(0x90), 0xBC] // U+897F <cjk>
	`誠`: [u8(0x90), 0xBD] // U+8AA0 <cjk>
	`誓`: [u8(0x90), 0xBE] // U+8A93 <cjk>
	`請`: [u8(0x90), 0xBF] // U+8ACB <cjk>
	`逝`: [u8(0x90), 0xC0] // U+901D <cjk>
	`醒`: [u8(0x90), 0xC1] // U+9192 <cjk>
	`青`: [u8(0x90), 0xC2] // U+9752 <cjk>
	`静`: [u8(0x90), 0xC3] // U+9759 <cjk>
	`斉`: [u8(0x90), 0xC4] // U+6589 <cjk>
	`税`: [u8(0x90), 0xC5] // U+7A0E <cjk>
	`脆`: [u8(0x90), 0xC6] // U+8106 <cjk>
	`隻`: [u8(0x90), 0xC7] // U+96BB <cjk>
	`席`: [u8(0x90), 0xC8] // U+5E2D <cjk>
	`惜`: [u8(0x90), 0xC9] // U+60DC <cjk>
	`戚`: [u8(0x90), 0xCA] // U+621A <cjk>
	`斥`: [u8(0x90), 0xCB] // U+65A5 <cjk>
	`昔`: [u8(0x90), 0xCC] // U+6614 <cjk>
	`析`: [u8(0x90), 0xCD] // U+6790 <cjk>
	`石`: [u8(0x90), 0xCE] // U+77F3 <cjk>
	`積`: [u8(0x90), 0xCF] // U+7A4D <cjk>
	`籍`: [u8(0x90), 0xD0] // U+7C4D <cjk>
	`績`: [u8(0x90), 0xD1] // U+7E3E <cjk>
	`脊`: [u8(0x90), 0xD2] // U+810A <cjk>
	`責`: [u8(0x90), 0xD3] // U+8CAC <cjk>
	`赤`: [u8(0x90), 0xD4] // U+8D64 <cjk>
	`跡`: [u8(0x90), 0xD5] // U+8DE1 <cjk>
	`蹟`: [u8(0x90), 0xD6] // U+8E5F <cjk>
	`碩`: [u8(0x90), 0xD7] // U+78A9 <cjk>
	`切`: [u8(0x90), 0xD8] // U+5207 <cjk>
	`拙`: [u8(0x90), 0xD9] // U+62D9 <cjk>
	`接`: [u8(0x90), 0xDA] // U+63A5 <cjk>
	`摂`: [u8(0x90), 0xDB] // U+6442 <cjk>
	`折`: [u8(0x90), 0xDC] // U+6298 <cjk>
	`設`: [u8(0x90), 0xDD] // U+8A2D <cjk>
	`窃`: [u8(0x90), 0xDE] // U+7A83 <cjk>
	`節`: [u8(0x90), 0xDF] // U+7BC0 <cjk>
	`説`: [u8(0x90), 0xE0] // U+8AAC <cjk>
	`雪`: [u8(0x90), 0xE1] // U+96EA <cjk>
	`絶`: [u8(0x90), 0xE2] // U+7D76 <cjk>
	`舌`: [u8(0x90), 0xE3] // U+820C <cjk>
	`蝉`: [u8(0x90), 0xE4] // U+8749 <cjk>
	`仙`: [u8(0x90), 0xE5] // U+4ED9 <cjk>
	`先`: [u8(0x90), 0xE6] // U+5148 <cjk>
	`千`: [u8(0x90), 0xE7] // U+5343 <cjk>
	`占`: [u8(0x90), 0xE8] // U+5360 <cjk>
	`宣`: [u8(0x90), 0xE9] // U+5BA3 <cjk>
	`専`: [u8(0x90), 0xEA] // U+5C02 <cjk>
	`尖`: [u8(0x90), 0xEB] // U+5C16 <cjk>
	`川`: [u8(0x90), 0xEC] // U+5DDD <cjk>
	`戦`: [u8(0x90), 0xED] // U+6226 <cjk>
	`扇`: [u8(0x90), 0xEE] // U+6247 <cjk>
	`撰`: [u8(0x90), 0xEF] // U+64B0 <cjk>
	`栓`: [u8(0x90), 0xF0] // U+6813 <cjk>
	`栴`: [u8(0x90), 0xF1] // U+6834 <cjk>
	`泉`: [u8(0x90), 0xF2] // U+6CC9 <cjk>
	`浅`: [u8(0x90), 0xF3] // U+6D45 <cjk>
	`洗`: [u8(0x90), 0xF4] // U+6D17 <cjk>
	`染`: [u8(0x90), 0xF5] // U+67D3 <cjk>
	`潜`: [u8(0x90), 0xF6] // U+6F5C <cjk>
	`煎`: [u8(0x90), 0xF7] // U+714E <cjk>
	`煽`: [u8(0x90), 0xF8] // U+717D <cjk>
	`旋`: [u8(0x90), 0xF9] // U+65CB <cjk>
	`穿`: [u8(0x90), 0xFA] // U+7A7F <cjk>
	`箭`: [u8(0x90), 0xFB] // U+7BAD <cjk>
	`線`: [u8(0x90), 0xFC] // U+7DDA <cjk>
	`繊`: [u8(0x91), 0x40] // U+7E4A <cjk>
	`羨`: [u8(0x91), 0x41] // U+7FA8 <cjk>
	`腺`: [u8(0x91), 0x42] // U+817A <cjk>
	`舛`: [u8(0x91), 0x43] // U+821B <cjk>
	`船`: [u8(0x91), 0x44] // U+8239 <cjk>
	`薦`: [u8(0x91), 0x45] // U+85A6 <cjk>
	`詮`: [u8(0x91), 0x46] // U+8A6E <cjk>
	`賎`: [u8(0x91), 0x47] // U+8CCE <cjk>
	`践`: [u8(0x91), 0x48] // U+8DF5 <cjk>
	`選`: [u8(0x91), 0x49] // U+9078 <cjk>
	`遷`: [u8(0x91), 0x4A] // U+9077 <cjk>
	`銭`: [u8(0x91), 0x4B] // U+92AD <cjk>
	`銑`: [u8(0x91), 0x4C] // U+9291 <cjk>
	`閃`: [u8(0x91), 0x4D] // U+9583 <cjk>
	`鮮`: [u8(0x91), 0x4E] // U+9BAE <cjk>
	`前`: [u8(0x91), 0x4F] // U+524D <cjk>
	`善`: [u8(0x91), 0x50] // U+5584 <cjk>
	`漸`: [u8(0x91), 0x51] // U+6F38 <cjk>
	`然`: [u8(0x91), 0x52] // U+7136 <cjk>
	`全`: [u8(0x91), 0x53] // U+5168 <cjk>
	`禅`: [u8(0x91), 0x54] // U+7985 <cjk>
	`繕`: [u8(0x91), 0x55] // U+7E55 <cjk>
	`膳`: [u8(0x91), 0x56] // U+81B3 <cjk>
	`糎`: [u8(0x91), 0x57] // U+7CCE <cjk>
	`噌`: [u8(0x91), 0x58] // U+564C <cjk>
	`塑`: [u8(0x91), 0x59] // U+5851 <cjk>
	`岨`: [u8(0x91), 0x5A] // U+5CA8 <cjk>
	`措`: [u8(0x91), 0x5B] // U+63AA <cjk>
	`曾`: [u8(0x91), 0x5C] // U+66FE <cjk>
	`曽`: [u8(0x91), 0x5D] // U+66FD <cjk>
	`楚`: [u8(0x91), 0x5E] // U+695A <cjk>
	`狙`: [u8(0x91), 0x5F] // U+72D9 <cjk>
	`疏`: [u8(0x91), 0x60] // U+758F <cjk>
	`疎`: [u8(0x91), 0x61] // U+758E <cjk>
	`礎`: [u8(0x91), 0x62] // U+790E <cjk>
	`祖`: [u8(0x91), 0x63] // U+7956 <cjk>
	`租`: [u8(0x91), 0x64] // U+79DF <cjk>
	`粗`: [u8(0x91), 0x65] // U+7C97 <cjk>
	`素`: [u8(0x91), 0x66] // U+7D20 <cjk>
	`組`: [u8(0x91), 0x67] // U+7D44 <cjk>
	`蘇`: [u8(0x91), 0x68] // U+8607 <cjk>
	`訴`: [u8(0x91), 0x69] // U+8A34 <cjk>
	`阻`: [u8(0x91), 0x6A] // U+963B <cjk>
	`遡`: [u8(0x91), 0x6B] // U+9061 <cjk>
	`鼠`: [u8(0x91), 0x6C] // U+9F20 <cjk>
	`僧`: [u8(0x91), 0x6D] // U+50E7 <cjk>
	`創`: [u8(0x91), 0x6E] // U+5275 <cjk>
	`双`: [u8(0x91), 0x6F] // U+53CC <cjk>
	`叢`: [u8(0x91), 0x70] // U+53E2 <cjk>
	`倉`: [u8(0x91), 0x71] // U+5009 <cjk>
	`喪`: [u8(0x91), 0x72] // U+55AA <cjk>
	`壮`: [u8(0x91), 0x73] // U+58EE <cjk>
	`奏`: [u8(0x91), 0x74] // U+594F <cjk>
	`爽`: [u8(0x91), 0x75] // U+723D <cjk>
	`宋`: [u8(0x91), 0x76] // U+5B8B <cjk>
	`層`: [u8(0x91), 0x77] // U+5C64 <cjk>
	`匝`: [u8(0x91), 0x78] // U+531D <cjk>
	`惣`: [u8(0x91), 0x79] // U+60E3 <cjk>
	`想`: [u8(0x91), 0x7A] // U+60F3 <cjk>
	`捜`: [u8(0x91), 0x7B] // U+635C <cjk>
	`掃`: [u8(0x91), 0x7C] // U+6383 <cjk>
	`挿`: [u8(0x91), 0x7D] // U+633F <cjk>
	`掻`: [u8(0x91), 0x7E] // U+63BB <cjk>
	`操`: [u8(0x91), 0x80] // U+64CD <cjk>
	`早`: [u8(0x91), 0x81] // U+65E9 <cjk>
	`曹`: [u8(0x91), 0x82] // U+66F9 <cjk>
	`巣`: [u8(0x91), 0x83] // U+5DE3 <cjk>
	`槍`: [u8(0x91), 0x84] // U+69CD <cjk>
	`槽`: [u8(0x91), 0x85] // U+69FD <cjk>
	`漕`: [u8(0x91), 0x86] // U+6F15 <cjk>
	`燥`: [u8(0x91), 0x87] // U+71E5 <cjk>
	`争`: [u8(0x91), 0x88] // U+4E89 <cjk>
	`痩`: [u8(0x91), 0x89] // U+75E9 <cjk>
	`相`: [u8(0x91), 0x8A] // U+76F8 <cjk>
	`窓`: [u8(0x91), 0x8B] // U+7A93 <cjk>
	`糟`: [u8(0x91), 0x8C] // U+7CDF <cjk>
	`総`: [u8(0x91), 0x8D] // U+7DCF <cjk>
	`綜`: [u8(0x91), 0x8E] // U+7D9C <cjk>
	`聡`: [u8(0x91), 0x8F] // U+8061 <cjk>
	`草`: [u8(0x91), 0x90] // U+8349 <cjk>
	`荘`: [u8(0x91), 0x91] // U+8358 <cjk>
	`葬`: [u8(0x91), 0x92] // U+846C <cjk>
	`蒼`: [u8(0x91), 0x93] // U+84BC <cjk>
	`藻`: [u8(0x91), 0x94] // U+85FB <cjk>
	`装`: [u8(0x91), 0x95] // U+88C5 <cjk>
	`走`: [u8(0x91), 0x96] // U+8D70 <cjk>
	`送`: [u8(0x91), 0x97] // U+9001 <cjk>
	`遭`: [u8(0x91), 0x98] // U+906D <cjk>
	`鎗`: [u8(0x91), 0x99] // U+9397 <cjk>
	`霜`: [u8(0x91), 0x9A] // U+971C <cjk>
	`騒`: [u8(0x91), 0x9B] // U+9A12 <cjk>
	`像`: [u8(0x91), 0x9C] // U+50CF <cjk>
	`増`: [u8(0x91), 0x9D] // U+5897 <cjk>
	`憎`: [u8(0x91), 0x9E] // U+618E <cjk>
	`臓`: [u8(0x91), 0x9F] // U+81D3 <cjk>
	`蔵`: [u8(0x91), 0xA0] // U+8535 <cjk>
	`贈`: [u8(0x91), 0xA1] // U+8D08 <cjk>
	`造`: [u8(0x91), 0xA2] // U+9020 <cjk>
	`促`: [u8(0x91), 0xA3] // U+4FC3 <cjk>
	`側`: [u8(0x91), 0xA4] // U+5074 <cjk>
	`則`: [u8(0x91), 0xA5] // U+5247 <cjk>
	`即`: [u8(0x91), 0xA6] // U+5373 <cjk>
	`息`: [u8(0x91), 0xA7] // U+606F <cjk>
	`捉`: [u8(0x91), 0xA8] // U+6349 <cjk>
	`束`: [u8(0x91), 0xA9] // U+675F <cjk>
	`測`: [u8(0x91), 0xAA] // U+6E2C <cjk>
	`足`: [u8(0x91), 0xAB] // U+8DB3 <cjk>
	`速`: [u8(0x91), 0xAC] // U+901F <cjk>
	`俗`: [u8(0x91), 0xAD] // U+4FD7 <cjk>
	`属`: [u8(0x91), 0xAE] // U+5C5E <cjk>
	`賊`: [u8(0x91), 0xAF] // U+8CCA <cjk>
	`族`: [u8(0x91), 0xB0] // U+65CF <cjk>
	`続`: [u8(0x91), 0xB1] // U+7D9A <cjk>
	`卒`: [u8(0x91), 0xB2] // U+5352 <cjk>
	`袖`: [u8(0x91), 0xB3] // U+8896 <cjk>
	`其`: [u8(0x91), 0xB4] // U+5176 <cjk>
	`揃`: [u8(0x91), 0xB5] // U+63C3 <cjk>
	`存`: [u8(0x91), 0xB6] // U+5B58 <cjk>
	`孫`: [u8(0x91), 0xB7] // U+5B6B <cjk>
	`尊`: [u8(0x91), 0xB8] // U+5C0A <cjk>
	`損`: [u8(0x91), 0xB9] // U+640D <cjk>
	`村`: [u8(0x91), 0xBA] // U+6751 <cjk>
	`遜`: [u8(0x91), 0xBB] // U+905C <cjk>
	`他`: [u8(0x91), 0xBC] // U+4ED6 <cjk>
	`多`: [u8(0x91), 0xBD] // U+591A <cjk>
	`太`: [u8(0x91), 0xBE] // U+592A <cjk>
	`汰`: [u8(0x91), 0xBF] // U+6C70 <cjk>
	`詑`: [u8(0x91), 0xC0] // U+8A51 <cjk>
	`唾`: [u8(0x91), 0xC1] // U+553E <cjk>
	`堕`: [u8(0x91), 0xC2] // U+5815 <cjk>
	`妥`: [u8(0x91), 0xC3] // U+59A5 <cjk>
	`惰`: [u8(0x91), 0xC4] // U+60F0 <cjk>
	`打`: [u8(0x91), 0xC5] // U+6253 <cjk>
	`柁`: [u8(0x91), 0xC6] // U+67C1 <cjk>
	`舵`: [u8(0x91), 0xC7] // U+8235 <cjk>
	`楕`: [u8(0x91), 0xC8] // U+6955 <cjk>
	`陀`: [u8(0x91), 0xC9] // U+9640 <cjk>
	`駄`: [u8(0x91), 0xCA] // U+99C4 <cjk>
	`騨`: [u8(0x91), 0xCB] // U+9A28 <cjk>
	`体`: [u8(0x91), 0xCC] // U+4F53 <cjk>
	`堆`: [u8(0x91), 0xCD] // U+5806 <cjk>
	`対`: [u8(0x91), 0xCE] // U+5BFE <cjk>
	`耐`: [u8(0x91), 0xCF] // U+8010 <cjk>
	`岱`: [u8(0x91), 0xD0] // U+5CB1 <cjk>
	`帯`: [u8(0x91), 0xD1] // U+5E2F <cjk>
	`待`: [u8(0x91), 0xD2] // U+5F85 <cjk>
	`怠`: [u8(0x91), 0xD3] // U+6020 <cjk>
	`態`: [u8(0x91), 0xD4] // U+614B <cjk>
	`戴`: [u8(0x91), 0xD5] // U+6234 <cjk>
	`替`: [u8(0x91), 0xD6] // U+66FF <cjk>
	`泰`: [u8(0x91), 0xD7] // U+6CF0 <cjk>
	`滞`: [u8(0x91), 0xD8] // U+6EDE <cjk>
	`胎`: [u8(0x91), 0xD9] // U+80CE <cjk>
	`腿`: [u8(0x91), 0xDA] // U+817F <cjk>
	`苔`: [u8(0x91), 0xDB] // U+82D4 <cjk>
	`袋`: [u8(0x91), 0xDC] // U+888B <cjk>
	`貸`: [u8(0x91), 0xDD] // U+8CB8 <cjk>
	`退`: [u8(0x91), 0xDE] // U+9000 <cjk>
	`逮`: [u8(0x91), 0xDF] // U+902E <cjk>
	`隊`: [u8(0x91), 0xE0] // U+968A <cjk>
	`黛`: [u8(0x91), 0xE1] // U+9EDB <cjk>
	`鯛`: [u8(0x91), 0xE2] // U+9BDB <cjk>
	`代`: [u8(0x91), 0xE3] // U+4EE3 <cjk>
	`台`: [u8(0x91), 0xE4] // U+53F0 <cjk>
	`大`: [u8(0x91), 0xE5] // U+5927 <cjk>
	`第`: [u8(0x91), 0xE6] // U+7B2C <cjk>
	`醍`: [u8(0x91), 0xE7] // U+918D <cjk>
	`題`: [u8(0x91), 0xE8] // U+984C <cjk>
	`鷹`: [u8(0x91), 0xE9] // U+9DF9 <cjk>
	`滝`: [u8(0x91), 0xEA] // U+6EDD <cjk>
	`瀧`: [u8(0x91), 0xEB] // U+7027 <cjk>
	`卓`: [u8(0x91), 0xEC] // U+5353 <cjk>
	`啄`: [u8(0x91), 0xED] // U+5544 <cjk>
	`宅`: [u8(0x91), 0xEE] // U+5B85 <cjk>
	`托`: [u8(0x91), 0xEF] // U+6258 <cjk>
	`択`: [u8(0x91), 0xF0] // U+629E <cjk>
	`拓`: [u8(0x91), 0xF1] // U+62D3 <cjk>
	`沢`: [u8(0x91), 0xF2] // U+6CA2 <cjk>
	`濯`: [u8(0x91), 0xF3] // U+6FEF <cjk>
	`琢`: [u8(0x91), 0xF4] // U+7422 <cjk>
	`託`: [u8(0x91), 0xF5] // U+8A17 <cjk>
	`鐸`: [u8(0x91), 0xF6] // U+9438 <cjk>
	`濁`: [u8(0x91), 0xF7] // U+6FC1 <cjk>
	`諾`: [u8(0x91), 0xF8] // U+8AFE <cjk>
	`茸`: [u8(0x91), 0xF9] // U+8338 <cjk>
	`凧`: [u8(0x91), 0xFA] // U+51E7 <cjk>
	`蛸`: [u8(0x91), 0xFB] // U+86F8 <cjk>
	`只`: [u8(0x91), 0xFC] // U+53EA <cjk>
	`叩`: [u8(0x92), 0x40] // U+53E9 <cjk>
	`但`: [u8(0x92), 0x41] // U+4F46 <cjk>
	`達`: [u8(0x92), 0x42] // U+9054 <cjk>
	`辰`: [u8(0x92), 0x43] // U+8FB0 <cjk>
	`奪`: [u8(0x92), 0x44] // U+596A <cjk>
	`脱`: [u8(0x92), 0x45] // U+8131 <cjk>
	`巽`: [u8(0x92), 0x46] // U+5DFD <cjk>
	`竪`: [u8(0x92), 0x47] // U+7AEA <cjk>
	`辿`: [u8(0x92), 0x48] // U+8FBF <cjk>
	`棚`: [u8(0x92), 0x49] // U+68DA <cjk>
	`谷`: [u8(0x92), 0x4A] // U+8C37 <cjk>
	`狸`: [u8(0x92), 0x4B] // U+72F8 <cjk>
	`鱈`: [u8(0x92), 0x4C] // U+9C48 <cjk>
	`樽`: [u8(0x92), 0x4D] // U+6A3D <cjk>
	`誰`: [u8(0x92), 0x4E] // U+8AB0 <cjk>
	`丹`: [u8(0x92), 0x4F] // U+4E39 <cjk>
	`単`: [u8(0x92), 0x50] // U+5358 <cjk>
	`嘆`: [u8(0x92), 0x51] // U+5606 <cjk>
	`坦`: [u8(0x92), 0x52] // U+5766 <cjk>
	`担`: [u8(0x92), 0x53] // U+62C5 <cjk>
	`探`: [u8(0x92), 0x54] // U+63A2 <cjk>
	`旦`: [u8(0x92), 0x55] // U+65E6 <cjk>
	`歎`: [u8(0x92), 0x56] // U+6B4E <cjk>
	`淡`: [u8(0x92), 0x57] // U+6DE1 <cjk>
	`湛`: [u8(0x92), 0x58] // U+6E5B <cjk>
	`炭`: [u8(0x92), 0x59] // U+70AD <cjk>
	`短`: [u8(0x92), 0x5A] // U+77ED <cjk>
	`端`: [u8(0x92), 0x5B] // U+7AEF <cjk>
	`箪`: [u8(0x92), 0x5C] // U+7BAA <cjk>
	`綻`: [u8(0x92), 0x5D] // U+7DBB <cjk>
	`耽`: [u8(0x92), 0x5E] // U+803D <cjk>
	`胆`: [u8(0x92), 0x5F] // U+80C6 <cjk>
	`蛋`: [u8(0x92), 0x60] // U+86CB <cjk>
	`誕`: [u8(0x92), 0x61] // U+8A95 <cjk>
	`鍛`: [u8(0x92), 0x62] // U+935B <cjk>
	`団`: [u8(0x92), 0x63] // U+56E3 <cjk>
	`壇`: [u8(0x92), 0x64] // U+58C7 <cjk>
	`弾`: [u8(0x92), 0x65] // U+5F3E <cjk>
	`断`: [u8(0x92), 0x66] // U+65AD <cjk>
	`暖`: [u8(0x92), 0x67] // U+6696 <cjk>
	`檀`: [u8(0x92), 0x68] // U+6A80 <cjk>
	`段`: [u8(0x92), 0x69] // U+6BB5 <cjk>
	`男`: [u8(0x92), 0x6A] // U+7537 <cjk>
	`談`: [u8(0x92), 0x6B] // U+8AC7 <cjk>
	`値`: [u8(0x92), 0x6C] // U+5024 <cjk>
	`知`: [u8(0x92), 0x6D] // U+77E5 <cjk>
	`地`: [u8(0x92), 0x6E] // U+5730 <cjk>
	`弛`: [u8(0x92), 0x6F] // U+5F1B <cjk>
	`恥`: [u8(0x92), 0x70] // U+6065 <cjk>
	`智`: [u8(0x92), 0x71] // U+667A <cjk>
	`池`: [u8(0x92), 0x72] // U+6C60 <cjk>
	`痴`: [u8(0x92), 0x73] // U+75F4 <cjk>
	`稚`: [u8(0x92), 0x74] // U+7A1A <cjk>
	`置`: [u8(0x92), 0x75] // U+7F6E <cjk>
	`致`: [u8(0x92), 0x76] // U+81F4 <cjk>
	`蜘`: [u8(0x92), 0x77] // U+8718 <cjk>
	`遅`: [u8(0x92), 0x78] // U+9045 <cjk>
	`馳`: [u8(0x92), 0x79] // U+99B3 <cjk>
	`築`: [u8(0x92), 0x7A] // U+7BC9 <cjk>
	`畜`: [u8(0x92), 0x7B] // U+755C <cjk>
	`竹`: [u8(0x92), 0x7C] // U+7AF9 <cjk>
	`筑`: [u8(0x92), 0x7D] // U+7B51 <cjk>
	`蓄`: [u8(0x92), 0x7E] // U+84C4 <cjk>
	`逐`: [u8(0x92), 0x80] // U+9010 <cjk>
	`秩`: [u8(0x92), 0x81] // U+79E9 <cjk>
	`窒`: [u8(0x92), 0x82] // U+7A92 <cjk>
	`茶`: [u8(0x92), 0x83] // U+8336 <cjk>
	`嫡`: [u8(0x92), 0x84] // U+5AE1 <cjk>
	`着`: [u8(0x92), 0x85] // U+7740 <cjk>
	`中`: [u8(0x92), 0x86] // U+4E2D <cjk>
	`仲`: [u8(0x92), 0x87] // U+4EF2 <cjk>
	`宙`: [u8(0x92), 0x88] // U+5B99 <cjk>
	`忠`: [u8(0x92), 0x89] // U+5FE0 <cjk>
	`抽`: [u8(0x92), 0x8A] // U+62BD <cjk>
	`昼`: [u8(0x92), 0x8B] // U+663C <cjk>
	`柱`: [u8(0x92), 0x8C] // U+67F1 <cjk>
	`注`: [u8(0x92), 0x8D] // U+6CE8 <cjk>
	`虫`: [u8(0x92), 0x8E] // U+866B <cjk>
	`衷`: [u8(0x92), 0x8F] // U+8877 <cjk>
	`註`: [u8(0x92), 0x90] // U+8A3B <cjk>
	`酎`: [u8(0x92), 0x91] // U+914E <cjk>
	`鋳`: [u8(0x92), 0x92] // U+92F3 <cjk>
	`駐`: [u8(0x92), 0x93] // U+99D0 <cjk>
	`樗`: [u8(0x92), 0x94] // U+6A17 <cjk>
	`瀦`: [u8(0x92), 0x95] // U+7026 <cjk>
	`猪`: [u8(0x92), 0x96] // U+732A <cjk>
	`苧`: [u8(0x92), 0x97] // U+82E7 <cjk>
	`著`: [u8(0x92), 0x98] // U+8457 <cjk>
	`貯`: [u8(0x92), 0x99] // U+8CAF <cjk>
	`丁`: [u8(0x92), 0x9A] // U+4E01 <cjk>
	`兆`: [u8(0x92), 0x9B] // U+5146 <cjk>
	`凋`: [u8(0x92), 0x9C] // U+51CB <cjk>
	`喋`: [u8(0x92), 0x9D] // U+558B <cjk>
	`寵`: [u8(0x92), 0x9E] // U+5BF5 <cjk>
	`帖`: [u8(0x92), 0x9F] // U+5E16 <cjk>
	`帳`: [u8(0x92), 0xA0] // U+5E33 <cjk>
	`庁`: [u8(0x92), 0xA1] // U+5E81 <cjk>
	`弔`: [u8(0x92), 0xA2] // U+5F14 <cjk>
	`張`: [u8(0x92), 0xA3] // U+5F35 <cjk>
	`彫`: [u8(0x92), 0xA4] // U+5F6B <cjk>
	`徴`: [u8(0x92), 0xA5] // U+5FB4 <cjk>
	`懲`: [u8(0x92), 0xA6] // U+61F2 <cjk>
	`挑`: [u8(0x92), 0xA7] // U+6311 <cjk>
	`暢`: [u8(0x92), 0xA8] // U+66A2 <cjk>
	`朝`: [u8(0x92), 0xA9] // U+671D <cjk>
	`潮`: [u8(0x92), 0xAA] // U+6F6E <cjk>
	`牒`: [u8(0x92), 0xAB] // U+7252 <cjk>
	`町`: [u8(0x92), 0xAC] // U+753A <cjk>
	`眺`: [u8(0x92), 0xAD] // U+773A <cjk>
	`聴`: [u8(0x92), 0xAE] // U+8074 <cjk>
	`脹`: [u8(0x92), 0xAF] // U+8139 <cjk>
	`腸`: [u8(0x92), 0xB0] // U+8178 <cjk>
	`蝶`: [u8(0x92), 0xB1] // U+8776 <cjk>
	`調`: [u8(0x92), 0xB2] // U+8ABF <cjk>
	`諜`: [u8(0x92), 0xB3] // U+8ADC <cjk>
	`超`: [u8(0x92), 0xB4] // U+8D85 <cjk>
	`跳`: [u8(0x92), 0xB5] // U+8DF3 <cjk>
	`銚`: [u8(0x92), 0xB6] // U+929A <cjk>
	`長`: [u8(0x92), 0xB7] // U+9577 <cjk>
	`頂`: [u8(0x92), 0xB8] // U+9802 <cjk>
	`鳥`: [u8(0x92), 0xB9] // U+9CE5 <cjk>
	`勅`: [u8(0x92), 0xBA] // U+52C5 <cjk>
	`捗`: [u8(0x92), 0xBB] // U+6357 <cjk>
	`直`: [u8(0x92), 0xBC] // U+76F4 <cjk>
	`朕`: [u8(0x92), 0xBD] // U+6715 <cjk>
	`沈`: [u8(0x92), 0xBE] // U+6C88 <cjk>
	`珍`: [u8(0x92), 0xBF] // U+73CD <cjk>
	`賃`: [u8(0x92), 0xC0] // U+8CC3 <cjk>
	`鎮`: [u8(0x92), 0xC1] // U+93AE <cjk>
	`陳`: [u8(0x92), 0xC2] // U+9673 <cjk>
	`津`: [u8(0x92), 0xC3] // U+6D25 <cjk>
	`墜`: [u8(0x92), 0xC4] // U+589C <cjk>
	`椎`: [u8(0x92), 0xC5] // U+690E <cjk>
	`槌`: [u8(0x92), 0xC6] // U+69CC <cjk>
	`追`: [u8(0x92), 0xC7] // U+8FFD <cjk>
	`鎚`: [u8(0x92), 0xC8] // U+939A <cjk>
	`痛`: [u8(0x92), 0xC9] // U+75DB <cjk>
	`通`: [u8(0x92), 0xCA] // U+901A <cjk>
	`塚`: [u8(0x92), 0xCB] // U+585A <cjk>
	`栂`: [u8(0x92), 0xCC] // U+6802 <cjk>
	`掴`: [u8(0x92), 0xCD] // U+63B4 <cjk>
	`槻`: [u8(0x92), 0xCE] // U+69FB <cjk>
	`佃`: [u8(0x92), 0xCF] // U+4F43 <cjk>
	`漬`: [u8(0x92), 0xD0] // U+6F2C <cjk>
	`柘`: [u8(0x92), 0xD1] // U+67D8 <cjk>
	`辻`: [u8(0x92), 0xD2] // U+8FBB <cjk>
	`蔦`: [u8(0x92), 0xD3] // U+8526 <cjk>
	`綴`: [u8(0x92), 0xD4] // U+7DB4 <cjk>
	`鍔`: [u8(0x92), 0xD5] // U+9354 <cjk>
	`椿`: [u8(0x92), 0xD6] // U+693F <cjk>
	`潰`: [u8(0x92), 0xD7] // U+6F70 <cjk>
	`坪`: [u8(0x92), 0xD8] // U+576A <cjk>
	`壷`: [u8(0x92), 0xD9] // U+58F7 <cjk>
	`嬬`: [u8(0x92), 0xDA] // U+5B2C <cjk>
	`紬`: [u8(0x92), 0xDB] // U+7D2C <cjk>
	`爪`: [u8(0x92), 0xDC] // U+722A <cjk>
	`吊`: [u8(0x92), 0xDD] // U+540A <cjk>
	`釣`: [u8(0x92), 0xDE] // U+91E3 <cjk>
	`鶴`: [u8(0x92), 0xDF] // U+9DB4 <cjk>
	`亭`: [u8(0x92), 0xE0] // U+4EAD <cjk>
	`低`: [u8(0x92), 0xE1] // U+4F4E <cjk>
	`停`: [u8(0x92), 0xE2] // U+505C <cjk>
	`偵`: [u8(0x92), 0xE3] // U+5075 <cjk>
	`剃`: [u8(0x92), 0xE4] // U+5243 <cjk>
	`貞`: [u8(0x92), 0xE5] // U+8C9E <cjk>
	`呈`: [u8(0x92), 0xE6] // U+5448 <cjk>
	`堤`: [u8(0x92), 0xE7] // U+5824 <cjk>
	`定`: [u8(0x92), 0xE8] // U+5B9A <cjk>
	`帝`: [u8(0x92), 0xE9] // U+5E1D <cjk>
	`底`: [u8(0x92), 0xEA] // U+5E95 <cjk>
	`庭`: [u8(0x92), 0xEB] // U+5EAD <cjk>
	`廷`: [u8(0x92), 0xEC] // U+5EF7 <cjk>
	`弟`: [u8(0x92), 0xED] // U+5F1F <cjk>
	`悌`: [u8(0x92), 0xEE] // U+608C <cjk>
	`抵`: [u8(0x92), 0xEF] // U+62B5 <cjk>
	`挺`: [u8(0x92), 0xF0] // U+633A <cjk>
	`提`: [u8(0x92), 0xF1] // U+63D0 <cjk>
	`梯`: [u8(0x92), 0xF2] // U+68AF <cjk>
	`汀`: [u8(0x92), 0xF3] // U+6C40 <cjk>
	`碇`: [u8(0x92), 0xF4] // U+7887 <cjk>
	`禎`: [u8(0x92), 0xF5] // U+798E <cjk>
	`程`: [u8(0x92), 0xF6] // U+7A0B <cjk>
	`締`: [u8(0x92), 0xF7] // U+7DE0 <cjk>
	`艇`: [u8(0x92), 0xF8] // U+8247 <cjk>
	`訂`: [u8(0x92), 0xF9] // U+8A02 <cjk>
	`諦`: [u8(0x92), 0xFA] // U+8AE6 <cjk>
	`蹄`: [u8(0x92), 0xFB] // U+8E44 <cjk>
	`逓`: [u8(0x92), 0xFC] // U+9013 <cjk>
	`邸`: [u8(0x93), 0x40] // U+90B8 <cjk>
	`鄭`: [u8(0x93), 0x41] // U+912D <cjk>
	`釘`: [u8(0x93), 0x42] // U+91D8 <cjk>
	`鼎`: [u8(0x93), 0x43] // U+9F0E <cjk>
	`泥`: [u8(0x93), 0x44] // U+6CE5 <cjk>
	`摘`: [u8(0x93), 0x45] // U+6458 <cjk>
	`擢`: [u8(0x93), 0x46] // U+64E2 <cjk>
	`敵`: [u8(0x93), 0x47] // U+6575 <cjk>
	`滴`: [u8(0x93), 0x48] // U+6EF4 <cjk>
	`的`: [u8(0x93), 0x49] // U+7684 <cjk>
	`笛`: [u8(0x93), 0x4A] // U+7B1B <cjk>
	`適`: [u8(0x93), 0x4B] // U+9069 <cjk>
	`鏑`: [u8(0x93), 0x4C] // U+93D1 <cjk>
	`溺`: [u8(0x93), 0x4D] // U+6EBA <cjk>
	`哲`: [u8(0x93), 0x4E] // U+54F2 <cjk>
	`徹`: [u8(0x93), 0x4F] // U+5FB9 <cjk>
	`撤`: [u8(0x93), 0x50] // U+64A4 <cjk>
	`轍`: [u8(0x93), 0x51] // U+8F4D <cjk>
	`迭`: [u8(0x93), 0x52] // U+8FED <cjk>
	`鉄`: [u8(0x93), 0x53] // U+9244 <cjk>
	`典`: [u8(0x93), 0x54] // U+5178 <cjk>
	`填`: [u8(0x93), 0x55] // U+586B <cjk>
	`天`: [u8(0x93), 0x56] // U+5929 <cjk>
	`展`: [u8(0x93), 0x57] // U+5C55 <cjk>
	`店`: [u8(0x93), 0x58] // U+5E97 <cjk>
	`添`: [u8(0x93), 0x59] // U+6DFB <cjk>
	`纏`: [u8(0x93), 0x5A] // U+7E8F <cjk>
	`甜`: [u8(0x93), 0x5B] // U+751C <cjk>
	`貼`: [u8(0x93), 0x5C] // U+8CBC <cjk>
	`転`: [u8(0x93), 0x5D] // U+8EE2 <cjk>
	`顛`: [u8(0x93), 0x5E] // U+985B <cjk>
	`点`: [u8(0x93), 0x5F] // U+70B9 <cjk>
	`伝`: [u8(0x93), 0x60] // U+4F1D <cjk>
	`殿`: [u8(0x93), 0x61] // U+6BBF <cjk>
	`澱`: [u8(0x93), 0x62] // U+6FB1 <cjk>
	`田`: [u8(0x93), 0x63] // U+7530 <cjk>
	`電`: [u8(0x93), 0x64] // U+96FB <cjk>
	`兎`: [u8(0x93), 0x65] // U+514E <cjk>
	`吐`: [u8(0x93), 0x66] // U+5410 <cjk>
	`堵`: [u8(0x93), 0x67] // U+5835 <cjk>
	`塗`: [u8(0x93), 0x68] // U+5857 <cjk>
	`妬`: [u8(0x93), 0x69] // U+59AC <cjk>
	`屠`: [u8(0x93), 0x6A] // U+5C60 <cjk>
	`徒`: [u8(0x93), 0x6B] // U+5F92 <cjk>
	`斗`: [u8(0x93), 0x6C] // U+6597 <cjk>
	`杜`: [u8(0x93), 0x6D] // U+675C <cjk>
	`渡`: [u8(0x93), 0x6E] // U+6E21 <cjk>
	`登`: [u8(0x93), 0x6F] // U+767B <cjk>
	`菟`: [u8(0x93), 0x70] // U+83DF <cjk>
	`賭`: [u8(0x93), 0x71] // U+8CED <cjk>
	`途`: [u8(0x93), 0x72] // U+9014 <cjk>
	`都`: [u8(0x93), 0x73] // U+90FD <cjk>
	`鍍`: [u8(0x93), 0x74] // U+934D <cjk>
	`砥`: [u8(0x93), 0x75] // U+7825 <cjk>
	`砺`: [u8(0x93), 0x76] // U+783A <cjk>
	`努`: [u8(0x93), 0x77] // U+52AA <cjk>
	`度`: [u8(0x93), 0x78] // U+5EA6 <cjk>
	`土`: [u8(0x93), 0x79] // U+571F <cjk>
	`奴`: [u8(0x93), 0x7A] // U+5974 <cjk>
	`怒`: [u8(0x93), 0x7B] // U+6012 <cjk>
	`倒`: [u8(0x93), 0x7C] // U+5012 <cjk>
	`党`: [u8(0x93), 0x7D] // U+515A <cjk>
	`冬`: [u8(0x93), 0x7E] // U+51AC <cjk>
	`凍`: [u8(0x93), 0x80] // U+51CD <cjk>
	`刀`: [u8(0x93), 0x81] // U+5200 <cjk>
	`唐`: [u8(0x93), 0x82] // U+5510 <cjk>
	`塔`: [u8(0x93), 0x83] // U+5854 <cjk>
	`塘`: [u8(0x93), 0x84] // U+5858 <cjk>
	`套`: [u8(0x93), 0x85] // U+5957 <cjk>
	`宕`: [u8(0x93), 0x86] // U+5B95 <cjk>
	`島`: [u8(0x93), 0x87] // U+5CF6 <cjk>
	`嶋`: [u8(0x93), 0x88] // U+5D8B <cjk>
	`悼`: [u8(0x93), 0x89] // U+60BC <cjk>
	`投`: [u8(0x93), 0x8A] // U+6295 <cjk>
	`搭`: [u8(0x93), 0x8B] // U+642D <cjk>
	`東`: [u8(0x93), 0x8C] // U+6771 <cjk>
	`桃`: [u8(0x93), 0x8D] // U+6843 <cjk>
	`梼`: [u8(0x93), 0x8E] // U+68BC <cjk>
	`棟`: [u8(0x93), 0x8F] // U+68DF <cjk>
	`盗`: [u8(0x93), 0x90] // U+76D7 <cjk>
	`淘`: [u8(0x93), 0x91] // U+6DD8 <cjk>
	`湯`: [u8(0x93), 0x92] // U+6E6F <cjk>
	`涛`: [u8(0x93), 0x93] // U+6D9B <cjk>
	`灯`: [u8(0x93), 0x94] // U+706F <cjk>
	`燈`: [u8(0x93), 0x95] // U+71C8 <cjk>
	`当`: [u8(0x93), 0x96] // U+5F53 <cjk>
	`痘`: [u8(0x93), 0x97] // U+75D8 <cjk>
	`祷`: [u8(0x93), 0x98] // U+7977 <cjk>
	`等`: [u8(0x93), 0x99] // U+7B49 <cjk>
	`答`: [u8(0x93), 0x9A] // U+7B54 <cjk>
	`筒`: [u8(0x93), 0x9B] // U+7B52 <cjk>
	`糖`: [u8(0x93), 0x9C] // U+7CD6 <cjk>
	`統`: [u8(0x93), 0x9D] // U+7D71 <cjk>
	`到`: [u8(0x93), 0x9E] // U+5230 <cjk>
	`董`: [u8(0x93), 0x9F] // U+8463 <cjk>
	`蕩`: [u8(0x93), 0xA0] // U+8569 <cjk>
	`藤`: [u8(0x93), 0xA1] // U+85E4 <cjk>
	`討`: [u8(0x93), 0xA2] // U+8A0E <cjk>
	`謄`: [u8(0x93), 0xA3] // U+8B04 <cjk>
	`豆`: [u8(0x93), 0xA4] // U+8C46 <cjk>
	`踏`: [u8(0x93), 0xA5] // U+8E0F <cjk>
	`逃`: [u8(0x93), 0xA6] // U+9003 <cjk>
	`透`: [u8(0x93), 0xA7] // U+900F <cjk>
	`鐙`: [u8(0x93), 0xA8] // U+9419 <cjk>
	`陶`: [u8(0x93), 0xA9] // U+9676 <cjk>
	`頭`: [u8(0x93), 0xAA] // U+982D <cjk>
	`騰`: [u8(0x93), 0xAB] // U+9A30 <cjk>
	`闘`: [u8(0x93), 0xAC] // U+95D8 <cjk>
	`働`: [u8(0x93), 0xAD] // U+50CD <cjk>
	`動`: [u8(0x93), 0xAE] // U+52D5 <cjk>
	`同`: [u8(0x93), 0xAF] // U+540C <cjk>
	`堂`: [u8(0x93), 0xB0] // U+5802 <cjk>
	`導`: [u8(0x93), 0xB1] // U+5C0E <cjk>
	`憧`: [u8(0x93), 0xB2] // U+61A7 <cjk>
	`撞`: [u8(0x93), 0xB3] // U+649E <cjk>
	`洞`: [u8(0x93), 0xB4] // U+6D1E <cjk>
	`瞳`: [u8(0x93), 0xB5] // U+77B3 <cjk>
	`童`: [u8(0x93), 0xB6] // U+7AE5 <cjk>
	`胴`: [u8(0x93), 0xB7] // U+80F4 <cjk>
	`萄`: [u8(0x93), 0xB8] // U+8404 <cjk>
	`道`: [u8(0x93), 0xB9] // U+9053 <cjk>
	`銅`: [u8(0x93), 0xBA] // U+9285 <cjk>
	`峠`: [u8(0x93), 0xBB] // U+5CE0 <cjk>
	`鴇`: [u8(0x93), 0xBC] // U+9D07 <cjk>
	`匿`: [u8(0x93), 0xBD] // U+533F <cjk>
	`得`: [u8(0x93), 0xBE] // U+5F97 <cjk>
	`徳`: [u8(0x93), 0xBF] // U+5FB3 <cjk>
	`涜`: [u8(0x93), 0xC0] // U+6D9C <cjk>
	`特`: [u8(0x93), 0xC1] // U+7279 <cjk>
	`督`: [u8(0x93), 0xC2] // U+7763 <cjk>
	`禿`: [u8(0x93), 0xC3] // U+79BF <cjk>
	`篤`: [u8(0x93), 0xC4] // U+7BE4 <cjk>
	`毒`: [u8(0x93), 0xC5] // U+6BD2 <cjk>
	`独`: [u8(0x93), 0xC6] // U+72EC <cjk>
	`読`: [u8(0x93), 0xC7] // U+8AAD <cjk>
	`栃`: [u8(0x93), 0xC8] // U+6803 <cjk>
	`橡`: [u8(0x93), 0xC9] // U+6A61 <cjk>
	`凸`: [u8(0x93), 0xCA] // U+51F8 <cjk>
	`突`: [u8(0x93), 0xCB] // U+7A81 <cjk>
	`椴`: [u8(0x93), 0xCC] // U+6934 <cjk>
	`届`: [u8(0x93), 0xCD] // U+5C4A <cjk>
	`鳶`: [u8(0x93), 0xCE] // U+9CF6 <cjk>
	`苫`: [u8(0x93), 0xCF] // U+82EB <cjk>
	`寅`: [u8(0x93), 0xD0] // U+5BC5 <cjk>
	`酉`: [u8(0x93), 0xD1] // U+9149 <cjk>
	`瀞`: [u8(0x93), 0xD2] // U+701E <cjk>
	`噸`: [u8(0x93), 0xD3] // U+5678 <cjk>
	`屯`: [u8(0x93), 0xD4] // U+5C6F <cjk>
	`惇`: [u8(0x93), 0xD5] // U+60C7 <cjk>
	`敦`: [u8(0x93), 0xD6] // U+6566 <cjk>
	`沌`: [u8(0x93), 0xD7] // U+6C8C <cjk>
	`豚`: [u8(0x93), 0xD8] // U+8C5A <cjk>
	`遁`: [u8(0x93), 0xD9] // U+9041 <cjk>
	`頓`: [u8(0x93), 0xDA] // U+9813 <cjk>
	`呑`: [u8(0x93), 0xDB] // U+5451 <cjk>
	`曇`: [u8(0x93), 0xDC] // U+66C7 <cjk>
	`鈍`: [u8(0x93), 0xDD] // U+920D <cjk>
	`奈`: [u8(0x93), 0xDE] // U+5948 <cjk>
	`那`: [u8(0x93), 0xDF] // U+90A3 <cjk>
	`内`: [u8(0x93), 0xE0] // U+5185 <cjk>
	`乍`: [u8(0x93), 0xE1] // U+4E4D <cjk>
	`凪`: [u8(0x93), 0xE2] // U+51EA <cjk>
	`薙`: [u8(0x93), 0xE3] // U+8599 <cjk>
	`謎`: [u8(0x93), 0xE4] // U+8B0E <cjk>
	`灘`: [u8(0x93), 0xE5] // U+7058 <cjk>
	`捺`: [u8(0x93), 0xE6] // U+637A <cjk>
	`鍋`: [u8(0x93), 0xE7] // U+934B <cjk>
	`楢`: [u8(0x93), 0xE8] // U+6962 <cjk>
	`馴`: [u8(0x93), 0xE9] // U+99B4 <cjk>
	`縄`: [u8(0x93), 0xEA] // U+7E04 <cjk>
	`畷`: [u8(0x93), 0xEB] // U+7577 <cjk>
	`南`: [u8(0x93), 0xEC] // U+5357 <cjk>
	`楠`: [u8(0x93), 0xED] // U+6960 <cjk>
	`軟`: [u8(0x93), 0xEE] // U+8EDF <cjk>
	`難`: [u8(0x93), 0xEF] // U+96E3 <cjk>
	`汝`: [u8(0x93), 0xF0] // U+6C5D <cjk>
	`二`: [u8(0x93), 0xF1] // U+4E8C <cjk>
	`尼`: [u8(0x93), 0xF2] // U+5C3C <cjk>
	`弐`: [u8(0x93), 0xF3] // U+5F10 <cjk>
	`迩`: [u8(0x93), 0xF4] // U+8FE9 <cjk>
	`匂`: [u8(0x93), 0xF5] // U+5302 <cjk>
	`賑`: [u8(0x93), 0xF6] // U+8CD1 <cjk>
	`肉`: [u8(0x93), 0xF7] // U+8089 <cjk>
	`虹`: [u8(0x93), 0xF8] // U+8679 <cjk>
	`廿`: [u8(0x93), 0xF9] // U+5EFF <cjk>
	`日`: [u8(0x93), 0xFA] // U+65E5 <cjk>
	`乳`: [u8(0x93), 0xFB] // U+4E73 <cjk>
	`入`: [u8(0x93), 0xFC] // U+5165 <cjk>
	`如`: [u8(0x94), 0x40] // U+5982 <cjk>
	`尿`: [u8(0x94), 0x41] // U+5C3F <cjk>
	`韮`: [u8(0x94), 0x42] // U+97EE <cjk>
	`任`: [u8(0x94), 0x43] // U+4EFB <cjk>
	`妊`: [u8(0x94), 0x44] // U+598A <cjk>
	`忍`: [u8(0x94), 0x45] // U+5FCD <cjk>
	`認`: [u8(0x94), 0x46] // U+8A8D <cjk>
	`濡`: [u8(0x94), 0x47] // U+6FE1 <cjk>
	`禰`: [u8(0x94), 0x48] // U+79B0 <cjk>
	`祢`: [u8(0x94), 0x49] // U+7962 <cjk>
	`寧`: [u8(0x94), 0x4A] // U+5BE7 <cjk>
	`葱`: [u8(0x94), 0x4B] // U+8471 <cjk>
	`猫`: [u8(0x94), 0x4C] // U+732B <cjk>
	`熱`: [u8(0x94), 0x4D] // U+71B1 <cjk>
	`年`: [u8(0x94), 0x4E] // U+5E74 <cjk>
	`念`: [u8(0x94), 0x4F] // U+5FF5 <cjk>
	`捻`: [u8(0x94), 0x50] // U+637B <cjk>
	`撚`: [u8(0x94), 0x51] // U+649A <cjk>
	`燃`: [u8(0x94), 0x52] // U+71C3 <cjk>
	`粘`: [u8(0x94), 0x53] // U+7C98 <cjk>
	`乃`: [u8(0x94), 0x54] // U+4E43 <cjk>
	`廼`: [u8(0x94), 0x55] // U+5EFC <cjk>
	`之`: [u8(0x94), 0x56] // U+4E4B <cjk>
	`埜`: [u8(0x94), 0x57] // U+57DC <cjk>
	`嚢`: [u8(0x94), 0x58] // U+56A2 <cjk>
	`悩`: [u8(0x94), 0x59] // U+60A9 <cjk>
	`濃`: [u8(0x94), 0x5A] // U+6FC3 <cjk>
	`納`: [u8(0x94), 0x5B] // U+7D0D <cjk>
	`能`: [u8(0x94), 0x5C] // U+80FD <cjk>
	`脳`: [u8(0x94), 0x5D] // U+8133 <cjk>
	`膿`: [u8(0x94), 0x5E] // U+81BF <cjk>
	`農`: [u8(0x94), 0x5F] // U+8FB2 <cjk>
	`覗`: [u8(0x94), 0x60] // U+8997 <cjk>
	`蚤`: [u8(0x94), 0x61] // U+86A4 <cjk>
	`巴`: [u8(0x94), 0x62] // U+5DF4 <cjk>
	`把`: [u8(0x94), 0x63] // U+628A <cjk>
	`播`: [u8(0x94), 0x64] // U+64AD <cjk>
	`覇`: [u8(0x94), 0x65] // U+8987 <cjk>
	`杷`: [u8(0x94), 0x66] // U+6777 <cjk>
	`波`: [u8(0x94), 0x67] // U+6CE2 <cjk>
	`派`: [u8(0x94), 0x68] // U+6D3E <cjk>
	`琶`: [u8(0x94), 0x69] // U+7436 <cjk>
	`破`: [u8(0x94), 0x6A] // U+7834 <cjk>
	`婆`: [u8(0x94), 0x6B] // U+5A46 <cjk>
	`罵`: [u8(0x94), 0x6C] // U+7F75 <cjk>
	`芭`: [u8(0x94), 0x6D] // U+82AD <cjk>
	`馬`: [u8(0x94), 0x6E] // U+99AC <cjk>
	`俳`: [u8(0x94), 0x6F] // U+4FF3 <cjk>
	`廃`: [u8(0x94), 0x70] // U+5EC3 <cjk>
	`拝`: [u8(0x94), 0x71] // U+62DD <cjk>
	`排`: [u8(0x94), 0x72] // U+6392 <cjk>
	`敗`: [u8(0x94), 0x73] // U+6557 <cjk>
	`杯`: [u8(0x94), 0x74] // U+676F <cjk>
	`盃`: [u8(0x94), 0x75] // U+76C3 <cjk>
	`牌`: [u8(0x94), 0x76] // U+724C <cjk>
	`背`: [u8(0x94), 0x77] // U+80CC <cjk>
	`肺`: [u8(0x94), 0x78] // U+80BA <cjk>
	`輩`: [u8(0x94), 0x79] // U+8F29 <cjk>
	`配`: [u8(0x94), 0x7A] // U+914D <cjk>
	`倍`: [u8(0x94), 0x7B] // U+500D <cjk>
	`培`: [u8(0x94), 0x7C] // U+57F9 <cjk>
	`媒`: [u8(0x94), 0x7D] // U+5A92 <cjk>
	`梅`: [u8(0x94), 0x7E] // U+6885 <cjk>
	`楳`: [u8(0x94), 0x80] // U+6973 <cjk>
	`煤`: [u8(0x94), 0x81] // U+7164 <cjk>
	`狽`: [u8(0x94), 0x82] // U+72FD <cjk>
	`買`: [u8(0x94), 0x83] // U+8CB7 <cjk>
	`売`: [u8(0x94), 0x84] // U+58F2 <cjk>
	`賠`: [u8(0x94), 0x85] // U+8CE0 <cjk>
	`陪`: [u8(0x94), 0x86] // U+966A <cjk>
	`這`: [u8(0x94), 0x87] // U+9019 <cjk>
	`蝿`: [u8(0x94), 0x88] // U+877F <cjk>
	`秤`: [u8(0x94), 0x89] // U+79E4 <cjk>
	`矧`: [u8(0x94), 0x8A] // U+77E7 <cjk>
	`萩`: [u8(0x94), 0x8B] // U+8429 <cjk>
	`伯`: [u8(0x94), 0x8C] // U+4F2F <cjk>
	`剥`: [u8(0x94), 0x8D] // U+5265 <cjk>
	`博`: [u8(0x94), 0x8E] // U+535A <cjk>
	`拍`: [u8(0x94), 0x8F] // U+62CD <cjk>
	`柏`: [u8(0x94), 0x90] // U+67CF <cjk>
	`泊`: [u8(0x94), 0x91] // U+6CCA <cjk>
	`白`: [u8(0x94), 0x92] // U+767D <cjk>
	`箔`: [u8(0x94), 0x93] // U+7B94 <cjk>
	`粕`: [u8(0x94), 0x94] // U+7C95 <cjk>
	`舶`: [u8(0x94), 0x95] // U+8236 <cjk>
	`薄`: [u8(0x94), 0x96] // U+8584 <cjk>
	`迫`: [u8(0x94), 0x97] // U+8FEB <cjk>
	`曝`: [u8(0x94), 0x98] // U+66DD <cjk>
	`漠`: [u8(0x94), 0x99] // U+6F20 <cjk>
	`爆`: [u8(0x94), 0x9A] // U+7206 <cjk>
	`縛`: [u8(0x94), 0x9B] // U+7E1B <cjk>
	`莫`: [u8(0x94), 0x9C] // U+83AB <cjk>
	`駁`: [u8(0x94), 0x9D] // U+99C1 <cjk>
	`麦`: [u8(0x94), 0x9E] // U+9EA6 <cjk>
	`函`: [u8(0x94), 0x9F] // U+51FD <cjk>
	`箱`: [u8(0x94), 0xA0] // U+7BB1 <cjk>
	`硲`: [u8(0x94), 0xA1] // U+7872 <cjk>
	`箸`: [u8(0x94), 0xA2] // U+7BB8 <cjk>
	`肇`: [u8(0x94), 0xA3] // U+8087 <cjk>
	`筈`: [u8(0x94), 0xA4] // U+7B48 <cjk>
	`櫨`: [u8(0x94), 0xA5] // U+6AE8 <cjk>
	`幡`: [u8(0x94), 0xA6] // U+5E61 <cjk>
	`肌`: [u8(0x94), 0xA7] // U+808C <cjk>
	`畑`: [u8(0x94), 0xA8] // U+7551 <cjk>
	`畠`: [u8(0x94), 0xA9] // U+7560 <cjk>
	`八`: [u8(0x94), 0xAA] // U+516B <cjk>
	`鉢`: [u8(0x94), 0xAB] // U+9262 <cjk>
	`溌`: [u8(0x94), 0xAC] // U+6E8C <cjk>
	`発`: [u8(0x94), 0xAD] // U+767A <cjk>
	`醗`: [u8(0x94), 0xAE] // U+9197 <cjk>
	`髪`: [u8(0x94), 0xAF] // U+9AEA <cjk>
	`伐`: [u8(0x94), 0xB0] // U+4F10 <cjk>
	`罰`: [u8(0x94), 0xB1] // U+7F70 <cjk>
	`抜`: [u8(0x94), 0xB2] // U+629C <cjk>
	`筏`: [u8(0x94), 0xB3] // U+7B4F <cjk>
	`閥`: [u8(0x94), 0xB4] // U+95A5 <cjk>
	`鳩`: [u8(0x94), 0xB5] // U+9CE9 <cjk>
	`噺`: [u8(0x94), 0xB6] // U+567A <cjk>
	`塙`: [u8(0x94), 0xB7] // U+5859 <cjk>
	`蛤`: [u8(0x94), 0xB8] // U+86E4 <cjk>
	`隼`: [u8(0x94), 0xB9] // U+96BC <cjk>
	`伴`: [u8(0x94), 0xBA] // U+4F34 <cjk>
	`判`: [u8(0x94), 0xBB] // U+5224 <cjk>
	`半`: [u8(0x94), 0xBC] // U+534A <cjk>
	`反`: [u8(0x94), 0xBD] // U+53CD <cjk>
	`叛`: [u8(0x94), 0xBE] // U+53DB <cjk>
	`帆`: [u8(0x94), 0xBF] // U+5E06 <cjk>
	`搬`: [u8(0x94), 0xC0] // U+642C <cjk>
	`斑`: [u8(0x94), 0xC1] // U+6591 <cjk>
	`板`: [u8(0x94), 0xC2] // U+677F <cjk>
	`氾`: [u8(0x94), 0xC3] // U+6C3E <cjk>
	`汎`: [u8(0x94), 0xC4] // U+6C4E <cjk>
	`版`: [u8(0x94), 0xC5] // U+7248 <cjk>
	`犯`: [u8(0x94), 0xC6] // U+72AF <cjk>
	`班`: [u8(0x94), 0xC7] // U+73ED <cjk>
	`畔`: [u8(0x94), 0xC8] // U+7554 <cjk>
	`繁`: [u8(0x94), 0xC9] // U+7E41 <cjk>
	`般`: [u8(0x94), 0xCA] // U+822C <cjk>
	`藩`: [u8(0x94), 0xCB] // U+85E9 <cjk>
	`販`: [u8(0x94), 0xCC] // U+8CA9 <cjk>
	`範`: [u8(0x94), 0xCD] // U+7BC4 <cjk>
	`釆`: [u8(0x94), 0xCE] // U+91C6 <cjk>
	`煩`: [u8(0x94), 0xCF] // U+7169 <cjk>
	`頒`: [u8(0x94), 0xD0] // U+9812 <cjk>
	`飯`: [u8(0x94), 0xD1] // U+98EF <cjk>
	`挽`: [u8(0x94), 0xD2] // U+633D <cjk>
	`晩`: [u8(0x94), 0xD3] // U+6669 <cjk>
	`番`: [u8(0x94), 0xD4] // U+756A <cjk>
	`盤`: [u8(0x94), 0xD5] // U+76E4 <cjk>
	`磐`: [u8(0x94), 0xD6] // U+78D0 <cjk>
	`蕃`: [u8(0x94), 0xD7] // U+8543 <cjk>
	`蛮`: [u8(0x94), 0xD8] // U+86EE <cjk>
	`匪`: [u8(0x94), 0xD9] // U+532A <cjk>
	`卑`: [u8(0x94), 0xDA] // U+5351 <cjk>
	`否`: [u8(0x94), 0xDB] // U+5426 <cjk>
	`妃`: [u8(0x94), 0xDC] // U+5983 <cjk>
	`庇`: [u8(0x94), 0xDD] // U+5E87 <cjk>
	`彼`: [u8(0x94), 0xDE] // U+5F7C <cjk>
	`悲`: [u8(0x94), 0xDF] // U+60B2 <cjk>
	`扉`: [u8(0x94), 0xE0] // U+6249 <cjk>
	`批`: [u8(0x94), 0xE1] // U+6279 <cjk>
	`披`: [u8(0x94), 0xE2] // U+62AB <cjk>
	`斐`: [u8(0x94), 0xE3] // U+6590 <cjk>
	`比`: [u8(0x94), 0xE4] // U+6BD4 <cjk>
	`泌`: [u8(0x94), 0xE5] // U+6CCC <cjk>
	`疲`: [u8(0x94), 0xE6] // U+75B2 <cjk>
	`皮`: [u8(0x94), 0xE7] // U+76AE <cjk>
	`碑`: [u8(0x94), 0xE8] // U+7891 <cjk>
	`秘`: [u8(0x94), 0xE9] // U+79D8 <cjk>
	`緋`: [u8(0x94), 0xEA] // U+7DCB <cjk>
	`罷`: [u8(0x94), 0xEB] // U+7F77 <cjk>
	`肥`: [u8(0x94), 0xEC] // U+80A5 <cjk>
	`被`: [u8(0x94), 0xED] // U+88AB <cjk>
	`誹`: [u8(0x94), 0xEE] // U+8AB9 <cjk>
	`費`: [u8(0x94), 0xEF] // U+8CBB <cjk>
	`避`: [u8(0x94), 0xF0] // U+907F <cjk>
	`非`: [u8(0x94), 0xF1] // U+975E <cjk>
	`飛`: [u8(0x94), 0xF2] // U+98DB <cjk>
	`樋`: [u8(0x94), 0xF3] // U+6A0B <cjk>
	`簸`: [u8(0x94), 0xF4] // U+7C38 <cjk>
	`備`: [u8(0x94), 0xF5] // U+5099 <cjk>
	`尾`: [u8(0x94), 0xF6] // U+5C3E <cjk>
	`微`: [u8(0x94), 0xF7] // U+5FAE <cjk>
	`枇`: [u8(0x94), 0xF8] // U+6787 <cjk>
	`毘`: [u8(0x94), 0xF9] // U+6BD8 <cjk>
	`琵`: [u8(0x94), 0xFA] // U+7435 <cjk>
	`眉`: [u8(0x94), 0xFB] // U+7709 <cjk>
	`美`: [u8(0x94), 0xFC] // U+7F8E <cjk>
	`鼻`: [u8(0x95), 0x40] // U+9F3B <cjk>
	`柊`: [u8(0x95), 0x41] // U+67CA <cjk>
	`稗`: [u8(0x95), 0x42] // U+7A17 <cjk>
	`匹`: [u8(0x95), 0x43] // U+5339 <cjk>
	`疋`: [u8(0x95), 0x44] // U+758B <cjk>
	`髭`: [u8(0x95), 0x45] // U+9AED <cjk>
	`彦`: [u8(0x95), 0x46] // U+5F66 <cjk>
	`膝`: [u8(0x95), 0x47] // U+819D <cjk>
	`菱`: [u8(0x95), 0x48] // U+83F1 <cjk>
	`肘`: [u8(0x95), 0x49] // U+8098 <cjk>
	`弼`: [u8(0x95), 0x4A] // U+5F3C <cjk>
	`必`: [u8(0x95), 0x4B] // U+5FC5 <cjk>
	`畢`: [u8(0x95), 0x4C] // U+7562 <cjk>
	`筆`: [u8(0x95), 0x4D] // U+7B46 <cjk>
	`逼`: [u8(0x95), 0x4E] // U+903C <cjk>
	`桧`: [u8(0x95), 0x4F] // U+6867 <cjk>
	`姫`: [u8(0x95), 0x50] // U+59EB <cjk>
	`媛`: [u8(0x95), 0x51] // U+5A9B <cjk>
	`紐`: [u8(0x95), 0x52] // U+7D10 <cjk>
	`百`: [u8(0x95), 0x53] // U+767E <cjk>
	`謬`: [u8(0x95), 0x54] // U+8B2C <cjk>
	`俵`: [u8(0x95), 0x55] // U+4FF5 <cjk>
	`彪`: [u8(0x95), 0x56] // U+5F6A <cjk>
	`標`: [u8(0x95), 0x57] // U+6A19 <cjk>
	`氷`: [u8(0x95), 0x58] // U+6C37 <cjk>
	`漂`: [u8(0x95), 0x59] // U+6F02 <cjk>
	`瓢`: [u8(0x95), 0x5A] // U+74E2 <cjk>
	`票`: [u8(0x95), 0x5B] // U+7968 <cjk>
	`表`: [u8(0x95), 0x5C] // U+8868 <cjk>
	`評`: [u8(0x95), 0x5D] // U+8A55 <cjk>
	`豹`: [u8(0x95), 0x5E] // U+8C79 <cjk>
	`廟`: [u8(0x95), 0x5F] // U+5EDF <cjk>
	`描`: [u8(0x95), 0x60] // U+63CF <cjk>
	`病`: [u8(0x95), 0x61] // U+75C5 <cjk>
	`秒`: [u8(0x95), 0x62] // U+79D2 <cjk>
	`苗`: [u8(0x95), 0x63] // U+82D7 <cjk>
	`錨`: [u8(0x95), 0x64] // U+9328 <cjk>
	`鋲`: [u8(0x95), 0x65] // U+92F2 <cjk>
	`蒜`: [u8(0x95), 0x66] // U+849C <cjk>
	`蛭`: [u8(0x95), 0x67] // U+86ED <cjk>
	`鰭`: [u8(0x95), 0x68] // U+9C2D <cjk>
	`品`: [u8(0x95), 0x69] // U+54C1 <cjk>
	`彬`: [u8(0x95), 0x6A] // U+5F6C <cjk>
	`斌`: [u8(0x95), 0x6B] // U+658C <cjk>
	`浜`: [u8(0x95), 0x6C] // U+6D5C <cjk>
	`瀕`: [u8(0x95), 0x6D] // U+7015 <cjk>
	`貧`: [u8(0x95), 0x6E] // U+8CA7 <cjk>
	`賓`: [u8(0x95), 0x6F] // U+8CD3 <cjk>
	`頻`: [u8(0x95), 0x70] // U+983B <cjk>
	`敏`: [u8(0x95), 0x71] // U+654F <cjk>
	`瓶`: [u8(0x95), 0x72] // U+74F6 <cjk>
	`不`: [u8(0x95), 0x73] // U+4E0D <cjk>
	`付`: [u8(0x95), 0x74] // U+4ED8 <cjk>
	`埠`: [u8(0x95), 0x75] // U+57E0 <cjk>
	`夫`: [u8(0x95), 0x76] // U+592B <cjk>
	`婦`: [u8(0x95), 0x77] // U+5A66 <cjk>
	`富`: [u8(0x95), 0x78] // U+5BCC <cjk>
	`冨`: [u8(0x95), 0x79] // U+51A8 <cjk>
	`布`: [u8(0x95), 0x7A] // U+5E03 <cjk>
	`府`: [u8(0x95), 0x7B] // U+5E9C <cjk>
	`怖`: [u8(0x95), 0x7C] // U+6016 <cjk>
	`扶`: [u8(0x95), 0x7D] // U+6276 <cjk>
	`敷`: [u8(0x95), 0x7E] // U+6577 <cjk>
	`斧`: [u8(0x95), 0x80] // U+65A7 <cjk>
	`普`: [u8(0x95), 0x81] // U+666E <cjk>
	`浮`: [u8(0x95), 0x82] // U+6D6E <cjk>
	`父`: [u8(0x95), 0x83] // U+7236 <cjk>
	`符`: [u8(0x95), 0x84] // U+7B26 <cjk>
	`腐`: [u8(0x95), 0x85] // U+8150 <cjk>
	`膚`: [u8(0x95), 0x86] // U+819A <cjk>
	`芙`: [u8(0x95), 0x87] // U+8299 <cjk>
	`譜`: [u8(0x95), 0x88] // U+8B5C <cjk>
	`負`: [u8(0x95), 0x89] // U+8CA0 <cjk>
	`賦`: [u8(0x95), 0x8A] // U+8CE6 <cjk>
	`赴`: [u8(0x95), 0x8B] // U+8D74 <cjk>
	`阜`: [u8(0x95), 0x8C] // U+961C <cjk>
	`附`: [u8(0x95), 0x8D] // U+9644 <cjk>
	`侮`: [u8(0x95), 0x8E] // U+4FAE <cjk>
	`撫`: [u8(0x95), 0x8F] // U+64AB <cjk>
	`武`: [u8(0x95), 0x90] // U+6B66 <cjk>
	`舞`: [u8(0x95), 0x91] // U+821E <cjk>
	`葡`: [u8(0x95), 0x92] // U+8461 <cjk>
	`蕪`: [u8(0x95), 0x93] // U+856A <cjk>
	`部`: [u8(0x95), 0x94] // U+90E8 <cjk>
	`封`: [u8(0x95), 0x95] // U+5C01 <cjk>
	`楓`: [u8(0x95), 0x96] // U+6953 <cjk>
	`風`: [u8(0x95), 0x97] // U+98A8 <cjk>
	`葺`: [u8(0x95), 0x98] // U+847A <cjk>
	`蕗`: [u8(0x95), 0x99] // U+8557 <cjk>
	`伏`: [u8(0x95), 0x9A] // U+4F0F <cjk>
	`副`: [u8(0x95), 0x9B] // U+526F <cjk>
	`復`: [u8(0x95), 0x9C] // U+5FA9 <cjk>
	`幅`: [u8(0x95), 0x9D] // U+5E45 <cjk>
	`服`: [u8(0x95), 0x9E] // U+670D <cjk>
	`福`: [u8(0x95), 0x9F] // U+798F <cjk>
	`腹`: [u8(0x95), 0xA0] // U+8179 <cjk>
	`複`: [u8(0x95), 0xA1] // U+8907 <cjk>
	`覆`: [u8(0x95), 0xA2] // U+8986 <cjk>
	`淵`: [u8(0x95), 0xA3] // U+6DF5 <cjk>
	`弗`: [u8(0x95), 0xA4] // U+5F17 <cjk>
	`払`: [u8(0x95), 0xA5] // U+6255 <cjk>
	`沸`: [u8(0x95), 0xA6] // U+6CB8 <cjk>
	`仏`: [u8(0x95), 0xA7] // U+4ECF <cjk>
	`物`: [u8(0x95), 0xA8] // U+7269 <cjk>
	`鮒`: [u8(0x95), 0xA9] // U+9B92 <cjk>
	`分`: [u8(0x95), 0xAA] // U+5206 <cjk>
	`吻`: [u8(0x95), 0xAB] // U+543B <cjk>
	`噴`: [u8(0x95), 0xAC] // U+5674 <cjk>
	`墳`: [u8(0x95), 0xAD] // U+58B3 <cjk>
	`憤`: [u8(0x95), 0xAE] // U+61A4 <cjk>
	`扮`: [u8(0x95), 0xAF] // U+626E <cjk>
	`焚`: [u8(0x95), 0xB0] // U+711A <cjk>
	`奮`: [u8(0x95), 0xB1] // U+596E <cjk>
	`粉`: [u8(0x95), 0xB2] // U+7C89 <cjk>
	`糞`: [u8(0x95), 0xB3] // U+7CDE <cjk>
	`紛`: [u8(0x95), 0xB4] // U+7D1B <cjk>
	`雰`: [u8(0x95), 0xB5] // U+96F0 <cjk>
	`文`: [u8(0x95), 0xB6] // U+6587 <cjk>
	`聞`: [u8(0x95), 0xB7] // U+805E <cjk>
	`丙`: [u8(0x95), 0xB8] // U+4E19 <cjk>
	`併`: [u8(0x95), 0xB9] // U+4F75 <cjk>
	`兵`: [u8(0x95), 0xBA] // U+5175 <cjk>
	`塀`: [u8(0x95), 0xBB] // U+5840 <cjk>
	`幣`: [u8(0x95), 0xBC] // U+5E63 <cjk>
	`平`: [u8(0x95), 0xBD] // U+5E73 <cjk>
	`弊`: [u8(0x95), 0xBE] // U+5F0A <cjk>
	`柄`: [u8(0x95), 0xBF] // U+67C4 <cjk>
	`並`: [u8(0x95), 0xC0] // U+4E26 <cjk>
	`蔽`: [u8(0x95), 0xC1] // U+853D <cjk>
	`閉`: [u8(0x95), 0xC2] // U+9589 <cjk>
	`陛`: [u8(0x95), 0xC3] // U+965B <cjk>
	`米`: [u8(0x95), 0xC4] // U+7C73 <cjk>
	`頁`: [u8(0x95), 0xC5] // U+9801 <cjk>
	`僻`: [u8(0x95), 0xC6] // U+50FB <cjk>
	`壁`: [u8(0x95), 0xC7] // U+58C1 <cjk>
	`癖`: [u8(0x95), 0xC8] // U+7656 <cjk>
	`碧`: [u8(0x95), 0xC9] // U+78A7 <cjk>
	`別`: [u8(0x95), 0xCA] // U+5225 <cjk>
	`瞥`: [u8(0x95), 0xCB] // U+77A5 <cjk>
	`蔑`: [u8(0x95), 0xCC] // U+8511 <cjk>
	`箆`: [u8(0x95), 0xCD] // U+7B86 <cjk>
	`偏`: [u8(0x95), 0xCE] // U+504F <cjk>
	`変`: [u8(0x95), 0xCF] // U+5909 <cjk>
	`片`: [u8(0x95), 0xD0] // U+7247 <cjk>
	`篇`: [u8(0x95), 0xD1] // U+7BC7 <cjk>
	`編`: [u8(0x95), 0xD2] // U+7DE8 <cjk>
	`辺`: [u8(0x95), 0xD3] // U+8FBA <cjk>
	`返`: [u8(0x95), 0xD4] // U+8FD4 <cjk>
	`遍`: [u8(0x95), 0xD5] // U+904D <cjk>
	`便`: [u8(0x95), 0xD6] // U+4FBF <cjk>
	`勉`: [u8(0x95), 0xD7] // U+52C9 <cjk>
	`娩`: [u8(0x95), 0xD8] // U+5A29 <cjk>
	`弁`: [u8(0x95), 0xD9] // U+5F01 <cjk>
	`鞭`: [u8(0x95), 0xDA] // U+97AD <cjk>
	`保`: [u8(0x95), 0xDB] // U+4FDD <cjk>
	`舗`: [u8(0x95), 0xDC] // U+8217 <cjk>
	`鋪`: [u8(0x95), 0xDD] // U+92EA <cjk>
	`圃`: [u8(0x95), 0xDE] // U+5703 <cjk>
	`捕`: [u8(0x95), 0xDF] // U+6355 <cjk>
	`歩`: [u8(0x95), 0xE0] // U+6B69 <cjk>
	`甫`: [u8(0x95), 0xE1] // U+752B <cjk>
	`補`: [u8(0x95), 0xE2] // U+88DC <cjk>
	`輔`: [u8(0x95), 0xE3] // U+8F14 <cjk>
	`穂`: [u8(0x95), 0xE4] // U+7A42 <cjk>
	`募`: [u8(0x95), 0xE5] // U+52DF <cjk>
	`墓`: [u8(0x95), 0xE6] // U+5893 <cjk>
	`慕`: [u8(0x95), 0xE7] // U+6155 <cjk>
	`戊`: [u8(0x95), 0xE8] // U+620A <cjk>
	`暮`: [u8(0x95), 0xE9] // U+66AE <cjk>
	`母`: [u8(0x95), 0xEA] // U+6BCD <cjk>
	`簿`: [u8(0x95), 0xEB] // U+7C3F <cjk>
	`菩`: [u8(0x95), 0xEC] // U+83E9 <cjk>
	`倣`: [u8(0x95), 0xED] // U+5023 <cjk>
	`俸`: [u8(0x95), 0xEE] // U+4FF8 <cjk>
	`包`: [u8(0x95), 0xEF] // U+5305 <cjk>
	`呆`: [u8(0x95), 0xF0] // U+5446 <cjk>
	`報`: [u8(0x95), 0xF1] // U+5831 <cjk>
	`奉`: [u8(0x95), 0xF2] // U+5949 <cjk>
	`宝`: [u8(0x95), 0xF3] // U+5B9D <cjk>
	`峰`: [u8(0x95), 0xF4] // U+5CF0 <cjk>
	`峯`: [u8(0x95), 0xF5] // U+5CEF <cjk>
	`崩`: [u8(0x95), 0xF6] // U+5D29 <cjk>
	`庖`: [u8(0x95), 0xF7] // U+5E96 <cjk>
	`抱`: [u8(0x95), 0xF8] // U+62B1 <cjk>
	`捧`: [u8(0x95), 0xF9] // U+6367 <cjk>
	`放`: [u8(0x95), 0xFA] // U+653E <cjk>
	`方`: [u8(0x95), 0xFB] // U+65B9 <cjk>
	`朋`: [u8(0x95), 0xFC] // U+670B <cjk>
	`法`: [u8(0x96), 0x40] // U+6CD5 <cjk>
	`泡`: [u8(0x96), 0x41] // U+6CE1 <cjk>
	`烹`: [u8(0x96), 0x42] // U+70F9 <cjk>
	`砲`: [u8(0x96), 0x43] // U+7832 <cjk>
	`縫`: [u8(0x96), 0x44] // U+7E2B <cjk>
	`胞`: [u8(0x96), 0x45] // U+80DE <cjk>
	`芳`: [u8(0x96), 0x46] // U+82B3 <cjk>
	`萌`: [u8(0x96), 0x47] // U+840C <cjk>
	`蓬`: [u8(0x96), 0x48] // U+84EC <cjk>
	`蜂`: [u8(0x96), 0x49] // U+8702 <cjk>
	`褒`: [u8(0x96), 0x4A] // U+8912 <cjk>
	`訪`: [u8(0x96), 0x4B] // U+8A2A <cjk>
	`豊`: [u8(0x96), 0x4C] // U+8C4A <cjk>
	`邦`: [u8(0x96), 0x4D] // U+90A6 <cjk>
	`鋒`: [u8(0x96), 0x4E] // U+92D2 <cjk>
	`飽`: [u8(0x96), 0x4F] // U+98FD <cjk>
	`鳳`: [u8(0x96), 0x50] // U+9CF3 <cjk>
	`鵬`: [u8(0x96), 0x51] // U+9D6C <cjk>
	`乏`: [u8(0x96), 0x52] // U+4E4F <cjk>
	`亡`: [u8(0x96), 0x53] // U+4EA1 <cjk>
	`傍`: [u8(0x96), 0x54] // U+508D <cjk>
	`剖`: [u8(0x96), 0x55] // U+5256 <cjk>
	`坊`: [u8(0x96), 0x56] // U+574A <cjk>
	`妨`: [u8(0x96), 0x57] // U+59A8 <cjk>
	`帽`: [u8(0x96), 0x58] // U+5E3D <cjk>
	`忘`: [u8(0x96), 0x59] // U+5FD8 <cjk>
	`忙`: [u8(0x96), 0x5A] // U+5FD9 <cjk>
	`房`: [u8(0x96), 0x5B] // U+623F <cjk>
	`暴`: [u8(0x96), 0x5C] // U+66B4 <cjk>
	`望`: [u8(0x96), 0x5D] // U+671B <cjk>
	`某`: [u8(0x96), 0x5E] // U+67D0 <cjk>
	`棒`: [u8(0x96), 0x5F] // U+68D2 <cjk>
	`冒`: [u8(0x96), 0x60] // U+5192 <cjk>
	`紡`: [u8(0x96), 0x61] // U+7D21 <cjk>
	`肪`: [u8(0x96), 0x62] // U+80AA <cjk>
	`膨`: [u8(0x96), 0x63] // U+81A8 <cjk>
	`謀`: [u8(0x96), 0x64] // U+8B00 <cjk>
	`貌`: [u8(0x96), 0x65] // U+8C8C <cjk>
	`貿`: [u8(0x96), 0x66] // U+8CBF <cjk>
	`鉾`: [u8(0x96), 0x67] // U+927E <cjk>
	`防`: [u8(0x96), 0x68] // U+9632 <cjk>
	`吠`: [u8(0x96), 0x69] // U+5420 <cjk>
	`頬`: [u8(0x96), 0x6A] // U+982C <cjk>
	`北`: [u8(0x96), 0x6B] // U+5317 <cjk>
	`僕`: [u8(0x96), 0x6C] // U+50D5 <cjk>
	`卜`: [u8(0x96), 0x6D] // U+535C <cjk>
	`墨`: [u8(0x96), 0x6E] // U+58A8 <cjk>
	`撲`: [u8(0x96), 0x6F] // U+64B2 <cjk>
	`朴`: [u8(0x96), 0x70] // U+6734 <cjk>
	`牧`: [u8(0x96), 0x71] // U+7267 <cjk>
	`睦`: [u8(0x96), 0x72] // U+7766 <cjk>
	`穆`: [u8(0x96), 0x73] // U+7A46 <cjk>
	`釦`: [u8(0x96), 0x74] // U+91E6 <cjk>
	`勃`: [u8(0x96), 0x75] // U+52C3 <cjk>
	`没`: [u8(0x96), 0x76] // U+6CA1 <cjk>
	`殆`: [u8(0x96), 0x77] // U+6B86 <cjk>
	`堀`: [u8(0x96), 0x78] // U+5800 <cjk>
	`幌`: [u8(0x96), 0x79] // U+5E4C <cjk>
	`奔`: [u8(0x96), 0x7A] // U+5954 <cjk>
	`本`: [u8(0x96), 0x7B] // U+672C <cjk>
	`翻`: [u8(0x96), 0x7C] // U+7FFB <cjk>
	`凡`: [u8(0x96), 0x7D] // U+51E1 <cjk>
	`盆`: [u8(0x96), 0x7E] // U+76C6 <cjk>
	`摩`: [u8(0x96), 0x80] // U+6469 <cjk>
	`磨`: [u8(0x96), 0x81] // U+78E8 <cjk>
	`魔`: [u8(0x96), 0x82] // U+9B54 <cjk>
	`麻`: [u8(0x96), 0x83] // U+9EBB <cjk>
	`埋`: [u8(0x96), 0x84] // U+57CB <cjk>
	`妹`: [u8(0x96), 0x85] // U+59B9 <cjk>
	`昧`: [u8(0x96), 0x86] // U+6627 <cjk>
	`枚`: [u8(0x96), 0x87] // U+679A <cjk>
	`毎`: [u8(0x96), 0x88] // U+6BCE <cjk>
	`哩`: [u8(0x96), 0x89] // U+54E9 <cjk>
	`槙`: [u8(0x96), 0x8A] // U+69D9 <cjk>
	`幕`: [u8(0x96), 0x8B] // U+5E55 <cjk>
	`膜`: [u8(0x96), 0x8C] // U+819C <cjk>
	`枕`: [u8(0x96), 0x8D] // U+6795 <cjk>
	`鮪`: [u8(0x96), 0x8E] // U+9BAA <cjk>
	`柾`: [u8(0x96), 0x8F] // U+67FE <cjk>
	`鱒`: [u8(0x96), 0x90] // U+9C52 <cjk>
	`桝`: [u8(0x96), 0x91] // U+685D <cjk>
	`亦`: [u8(0x96), 0x92] // U+4EA6 <cjk>
	`俣`: [u8(0x96), 0x93] // U+4FE3 <cjk>
	`又`: [u8(0x96), 0x94] // U+53C8 <cjk>
	`抹`: [u8(0x96), 0x95] // U+62B9 <cjk>
	`末`: [u8(0x96), 0x96] // U+672B <cjk>
	`沫`: [u8(0x96), 0x97] // U+6CAB <cjk>
	`迄`: [u8(0x96), 0x98] // U+8FC4 <cjk>
	`侭`: [u8(0x96), 0x99] // U+4FAD <cjk>
	`繭`: [u8(0x96), 0x9A] // U+7E6D <cjk>
	`麿`: [u8(0x96), 0x9B] // U+9EBF <cjk>
	`万`: [u8(0x96), 0x9C] // U+4E07 <cjk>
	`慢`: [u8(0x96), 0x9D] // U+6162 <cjk>
	`満`: [u8(0x96), 0x9E] // U+6E80 <cjk>
	`漫`: [u8(0x96), 0x9F] // U+6F2B <cjk>
	`蔓`: [u8(0x96), 0xA0] // U+8513 <cjk>
	`味`: [u8(0x96), 0xA1] // U+5473 <cjk>
	`未`: [u8(0x96), 0xA2] // U+672A <cjk>
	`魅`: [u8(0x96), 0xA3] // U+9B45 <cjk>
	`巳`: [u8(0x96), 0xA4] // U+5DF3 <cjk>
	`箕`: [u8(0x96), 0xA5] // U+7B95 <cjk>
	`岬`: [u8(0x96), 0xA6] // U+5CAC <cjk>
	`密`: [u8(0x96), 0xA7] // U+5BC6 <cjk>
	`蜜`: [u8(0x96), 0xA8] // U+871C <cjk>
	`湊`: [u8(0x96), 0xA9] // U+6E4A <cjk>
	`蓑`: [u8(0x96), 0xAA] // U+84D1 <cjk>
	`稔`: [u8(0x96), 0xAB] // U+7A14 <cjk>
	`脈`: [u8(0x96), 0xAC] // U+8108 <cjk>
	`妙`: [u8(0x96), 0xAD] // U+5999 <cjk>
	`粍`: [u8(0x96), 0xAE] // U+7C8D <cjk>
	`民`: [u8(0x96), 0xAF] // U+6C11 <cjk>
	`眠`: [u8(0x96), 0xB0] // U+7720 <cjk>
	`務`: [u8(0x96), 0xB1] // U+52D9 <cjk>
	`夢`: [u8(0x96), 0xB2] // U+5922 <cjk>
	`無`: [u8(0x96), 0xB3] // U+7121 <cjk>
	`牟`: [u8(0x96), 0xB4] // U+725F <cjk>
	`矛`: [u8(0x96), 0xB5] // U+77DB <cjk>
	`霧`: [u8(0x96), 0xB6] // U+9727 <cjk>
	`鵡`: [u8(0x96), 0xB7] // U+9D61 <cjk>
	`椋`: [u8(0x96), 0xB8] // U+690B <cjk>
	`婿`: [u8(0x96), 0xB9] // U+5A7F <cjk>
	`娘`: [u8(0x96), 0xBA] // U+5A18 <cjk>
	`冥`: [u8(0x96), 0xBB] // U+51A5 <cjk>
	`名`: [u8(0x96), 0xBC] // U+540D <cjk>
	`命`: [u8(0x96), 0xBD] // U+547D <cjk>
	`明`: [u8(0x96), 0xBE] // U+660E <cjk>
	`盟`: [u8(0x96), 0xBF] // U+76DF <cjk>
	`迷`: [u8(0x96), 0xC0] // U+8FF7 <cjk>
	`銘`: [u8(0x96), 0xC1] // U+9298 <cjk>
	`鳴`: [u8(0x96), 0xC2] // U+9CF4 <cjk>
	`姪`: [u8(0x96), 0xC3] // U+59EA <cjk>
	`牝`: [u8(0x96), 0xC4] // U+725D <cjk>
	`滅`: [u8(0x96), 0xC5] // U+6EC5 <cjk>
	`免`: [u8(0x96), 0xC6] // U+514D <cjk>
	`棉`: [u8(0x96), 0xC7] // U+68C9 <cjk>
	`綿`: [u8(0x96), 0xC8] // U+7DBF <cjk>
	`緬`: [u8(0x96), 0xC9] // U+7DEC <cjk>
	`面`: [u8(0x96), 0xCA] // U+9762 <cjk>
	`麺`: [u8(0x96), 0xCB] // U+9EBA <cjk>
	`摸`: [u8(0x96), 0xCC] // U+6478 <cjk>
	`模`: [u8(0x96), 0xCD] // U+6A21 <cjk>
	`茂`: [u8(0x96), 0xCE] // U+8302 <cjk>
	`妄`: [u8(0x96), 0xCF] // U+5984 <cjk>
	`孟`: [u8(0x96), 0xD0] // U+5B5F <cjk>
	`毛`: [u8(0x96), 0xD1] // U+6BDB <cjk>
	`猛`: [u8(0x96), 0xD2] // U+731B <cjk>
	`盲`: [u8(0x96), 0xD3] // U+76F2 <cjk>
	`網`: [u8(0x96), 0xD4] // U+7DB2 <cjk>
	`耗`: [u8(0x96), 0xD5] // U+8017 <cjk>
	`蒙`: [u8(0x96), 0xD6] // U+8499 <cjk>
	`儲`: [u8(0x96), 0xD7] // U+5132 <cjk>
	`木`: [u8(0x96), 0xD8] // U+6728 <cjk>
	`黙`: [u8(0x96), 0xD9] // U+9ED9 <cjk>
	`目`: [u8(0x96), 0xDA] // U+76EE <cjk>
	`杢`: [u8(0x96), 0xDB] // U+6762 <cjk>
	`勿`: [u8(0x96), 0xDC] // U+52FF <cjk>
	`餅`: [u8(0x96), 0xDD] // U+9905 <cjk>
	`尤`: [u8(0x96), 0xDE] // U+5C24 <cjk>
	`戻`: [u8(0x96), 0xDF] // U+623B <cjk>
	`籾`: [u8(0x96), 0xE0] // U+7C7E <cjk>
	`貰`: [u8(0x96), 0xE1] // U+8CB0 <cjk>
	`問`: [u8(0x96), 0xE2] // U+554F <cjk>
	`悶`: [u8(0x96), 0xE3] // U+60B6 <cjk>
	`紋`: [u8(0x96), 0xE4] // U+7D0B <cjk>
	`門`: [u8(0x96), 0xE5] // U+9580 <cjk>
	`匁`: [u8(0x96), 0xE6] // U+5301 <cjk>
	`也`: [u8(0x96), 0xE7] // U+4E5F <cjk>
	`冶`: [u8(0x96), 0xE8] // U+51B6 <cjk>
	`夜`: [u8(0x96), 0xE9] // U+591C <cjk>
	`爺`: [u8(0x96), 0xEA] // U+723A <cjk>
	`耶`: [u8(0x96), 0xEB] // U+8036 <cjk>
	`野`: [u8(0x96), 0xEC] // U+91CE <cjk>
	`弥`: [u8(0x96), 0xED] // U+5F25 <cjk>
	`矢`: [u8(0x96), 0xEE] // U+77E2 <cjk>
	`厄`: [u8(0x96), 0xEF] // U+5384 <cjk>
	`役`: [u8(0x96), 0xF0] // U+5F79 <cjk>
	`約`: [u8(0x96), 0xF1] // U+7D04 <cjk>
	`薬`: [u8(0x96), 0xF2] // U+85AC <cjk>
	`訳`: [u8(0x96), 0xF3] // U+8A33 <cjk>
	`躍`: [u8(0x96), 0xF4] // U+8E8D <cjk>
	`靖`: [u8(0x96), 0xF5] // U+9756 <cjk>
	`柳`: [u8(0x96), 0xF6] // U+67F3 <cjk>
	`薮`: [u8(0x96), 0xF7] // U+85AE <cjk>
	`鑓`: [u8(0x96), 0xF8] // U+9453 <cjk>
	`愉`: [u8(0x96), 0xF9] // U+6109 <cjk>
	`愈`: [u8(0x96), 0xFA] // U+6108 <cjk>
	`油`: [u8(0x96), 0xFB] // U+6CB9 <cjk>
	`癒`: [u8(0x96), 0xFC] // U+7652 <cjk>
	`諭`: [u8(0x97), 0x40] // U+8AED <cjk>
	`輸`: [u8(0x97), 0x41] // U+8F38 <cjk>
	`唯`: [u8(0x97), 0x42] // U+552F <cjk>
	`佑`: [u8(0x97), 0x43] // U+4F51 <cjk>
	`優`: [u8(0x97), 0x44] // U+512A <cjk>
	`勇`: [u8(0x97), 0x45] // U+52C7 <cjk>
	`友`: [u8(0x97), 0x46] // U+53CB <cjk>
	`宥`: [u8(0x97), 0x47] // U+5BA5 <cjk>
	`幽`: [u8(0x97), 0x48] // U+5E7D <cjk>
	`悠`: [u8(0x97), 0x49] // U+60A0 <cjk>
	`憂`: [u8(0x97), 0x4A] // U+6182 <cjk>
	`揖`: [u8(0x97), 0x4B] // U+63D6 <cjk>
	`有`: [u8(0x97), 0x4C] // U+6709 <cjk>
	`柚`: [u8(0x97), 0x4D] // U+67DA <cjk>
	`湧`: [u8(0x97), 0x4E] // U+6E67 <cjk>
	`涌`: [u8(0x97), 0x4F] // U+6D8C <cjk>
	`猶`: [u8(0x97), 0x50] // U+7336 <cjk>
	`猷`: [u8(0x97), 0x51] // U+7337 <cjk>
	`由`: [u8(0x97), 0x52] // U+7531 <cjk>
	`祐`: [u8(0x97), 0x53] // U+7950 <cjk>
	`裕`: [u8(0x97), 0x54] // U+88D5 <cjk>
	`誘`: [u8(0x97), 0x55] // U+8A98 <cjk>
	`遊`: [u8(0x97), 0x56] // U+904A <cjk>
	`邑`: [u8(0x97), 0x57] // U+9091 <cjk>
	`郵`: [u8(0x97), 0x58] // U+90F5 <cjk>
	`雄`: [u8(0x97), 0x59] // U+96C4 <cjk>
	`融`: [u8(0x97), 0x5A] // U+878D <cjk>
	`夕`: [u8(0x97), 0x5B] // U+5915 <cjk>
	`予`: [u8(0x97), 0x5C] // U+4E88 <cjk>
	`余`: [u8(0x97), 0x5D] // U+4F59 <cjk>
	`与`: [u8(0x97), 0x5E] // U+4E0E <cjk>
	`誉`: [u8(0x97), 0x5F] // U+8A89 <cjk>
	`輿`: [u8(0x97), 0x60] // U+8F3F <cjk>
	`預`: [u8(0x97), 0x61] // U+9810 <cjk>
	`傭`: [u8(0x97), 0x62] // U+50AD <cjk>
	`幼`: [u8(0x97), 0x63] // U+5E7C <cjk>
	`妖`: [u8(0x97), 0x64] // U+5996 <cjk>
	`容`: [u8(0x97), 0x65] // U+5BB9 <cjk>
	`庸`: [u8(0x97), 0x66] // U+5EB8 <cjk>
	`揚`: [u8(0x97), 0x67] // U+63DA <cjk>
	`揺`: [u8(0x97), 0x68] // U+63FA <cjk>
	`擁`: [u8(0x97), 0x69] // U+64C1 <cjk>
	`曜`: [u8(0x97), 0x6A] // U+66DC <cjk>
	`楊`: [u8(0x97), 0x6B] // U+694A <cjk>
	`様`: [u8(0x97), 0x6C] // U+69D8 <cjk>
	`洋`: [u8(0x97), 0x6D] // U+6D0B <cjk>
	`溶`: [u8(0x97), 0x6E] // U+6EB6 <cjk>
	`熔`: [u8(0x97), 0x6F] // U+7194 <cjk>
	`用`: [u8(0x97), 0x70] // U+7528 <cjk>
	`窯`: [u8(0x97), 0x71] // U+7AAF <cjk>
	`羊`: [u8(0x97), 0x72] // U+7F8A <cjk>
	`耀`: [u8(0x97), 0x73] // U+8000 <cjk>
	`葉`: [u8(0x97), 0x74] // U+8449 <cjk>
	`蓉`: [u8(0x97), 0x75] // U+84C9 <cjk>
	`要`: [u8(0x97), 0x76] // U+8981 <cjk>
	`謡`: [u8(0x97), 0x77] // U+8B21 <cjk>
	`踊`: [u8(0x97), 0x78] // U+8E0A <cjk>
	`遥`: [u8(0x97), 0x79] // U+9065 <cjk>
	`陽`: [u8(0x97), 0x7A] // U+967D <cjk>
	`養`: [u8(0x97), 0x7B] // U+990A <cjk>
	`慾`: [u8(0x97), 0x7C] // U+617E <cjk>
	`抑`: [u8(0x97), 0x7D] // U+6291 <cjk>
	`欲`: [u8(0x97), 0x7E] // U+6B32 <cjk>
	`沃`: [u8(0x97), 0x80] // U+6C83 <cjk>
	`浴`: [u8(0x97), 0x81] // U+6D74 <cjk>
	`翌`: [u8(0x97), 0x82] // U+7FCC <cjk>
	`翼`: [u8(0x97), 0x83] // U+7FFC <cjk>
	`淀`: [u8(0x97), 0x84] // U+6DC0 <cjk>
	`羅`: [u8(0x97), 0x85] // U+7F85 <cjk>
	`螺`: [u8(0x97), 0x86] // U+87BA <cjk>
	`裸`: [u8(0x97), 0x87] // U+88F8 <cjk>
	`来`: [u8(0x97), 0x88] // U+6765 <cjk>
	`莱`: [u8(0x97), 0x89] // U+83B1 <cjk>
	`頼`: [u8(0x97), 0x8A] // U+983C <cjk>
	`雷`: [u8(0x97), 0x8B] // U+96F7 <cjk>
	`洛`: [u8(0x97), 0x8C] // U+6D1B <cjk>
	`絡`: [u8(0x97), 0x8D] // U+7D61 <cjk>
	`落`: [u8(0x97), 0x8E] // U+843D <cjk>
	`酪`: [u8(0x97), 0x8F] // U+916A <cjk>
	`乱`: [u8(0x97), 0x90] // U+4E71 <cjk>
	`卵`: [u8(0x97), 0x91] // U+5375 <cjk>
	`嵐`: [u8(0x97), 0x92] // U+5D50 <cjk>
	`欄`: [u8(0x97), 0x93] // U+6B04 <cjk>
	`濫`: [u8(0x97), 0x94] // U+6FEB <cjk>
	`藍`: [u8(0x97), 0x95] // U+85CD <cjk>
	`蘭`: [u8(0x97), 0x96] // U+862D <cjk>
	`覧`: [u8(0x97), 0x97] // U+89A7 <cjk>
	`利`: [u8(0x97), 0x98] // U+5229 <cjk>
	`吏`: [u8(0x97), 0x99] // U+540F <cjk>
	`履`: [u8(0x97), 0x9A] // U+5C65 <cjk>
	`李`: [u8(0x97), 0x9B] // U+674E <cjk>
	`梨`: [u8(0x97), 0x9C] // U+68A8 <cjk>
	`理`: [u8(0x97), 0x9D] // U+7406 <cjk>
	`璃`: [u8(0x97), 0x9E] // U+7483 <cjk>
	`痢`: [u8(0x97), 0x9F] // U+75E2 <cjk>
	`裏`: [u8(0x97), 0xA0] // U+88CF <cjk>
	`裡`: [u8(0x97), 0xA1] // U+88E1 <cjk>
	`里`: [u8(0x97), 0xA2] // U+91CC <cjk>
	`離`: [u8(0x97), 0xA3] // U+96E2 <cjk>
	`陸`: [u8(0x97), 0xA4] // U+9678 <cjk>
	`律`: [u8(0x97), 0xA5] // U+5F8B <cjk>
	`率`: [u8(0x97), 0xA6] // U+7387 <cjk>
	`立`: [u8(0x97), 0xA7] // U+7ACB <cjk>
	`葎`: [u8(0x97), 0xA8] // U+844E <cjk>
	`掠`: [u8(0x97), 0xA9] // U+63A0 <cjk>
	`略`: [u8(0x97), 0xAA] // U+7565 <cjk>
	`劉`: [u8(0x97), 0xAB] // U+5289 <cjk>
	`流`: [u8(0x97), 0xAC] // U+6D41 <cjk>
	`溜`: [u8(0x97), 0xAD] // U+6E9C <cjk>
	`琉`: [u8(0x97), 0xAE] // U+7409 <cjk>
	`留`: [u8(0x97), 0xAF] // U+7559 <cjk>
	`硫`: [u8(0x97), 0xB0] // U+786B <cjk>
	`粒`: [u8(0x97), 0xB1] // U+7C92 <cjk>
	`隆`: [u8(0x97), 0xB2] // U+9686 <cjk>
	`竜`: [u8(0x97), 0xB3] // U+7ADC <cjk>
	`龍`: [u8(0x97), 0xB4] // U+9F8D <cjk>
	`侶`: [u8(0x97), 0xB5] // U+4FB6 <cjk>
	`慮`: [u8(0x97), 0xB6] // U+616E <cjk>
	`旅`: [u8(0x97), 0xB7] // U+65C5 <cjk>
	`虜`: [u8(0x97), 0xB8] // U+865C <cjk>
	`了`: [u8(0x97), 0xB9] // U+4E86 <cjk>
	`亮`: [u8(0x97), 0xBA] // U+4EAE <cjk>
	`僚`: [u8(0x97), 0xBB] // U+50DA <cjk>
	`両`: [u8(0x97), 0xBC] // U+4E21 <cjk>
	`凌`: [u8(0x97), 0xBD] // U+51CC <cjk>
	`寮`: [u8(0x97), 0xBE] // U+5BEE <cjk>
	`料`: [u8(0x97), 0xBF] // U+6599 <cjk>
	`梁`: [u8(0x97), 0xC0] // U+6881 <cjk>
	`涼`: [u8(0x97), 0xC1] // U+6DBC <cjk>
	`猟`: [u8(0x97), 0xC2] // U+731F <cjk>
	`療`: [u8(0x97), 0xC3] // U+7642 <cjk>
	`瞭`: [u8(0x97), 0xC4] // U+77AD <cjk>
	`稜`: [u8(0x97), 0xC5] // U+7A1C <cjk>
	`糧`: [u8(0x97), 0xC6] // U+7CE7 <cjk>
	`良`: [u8(0x97), 0xC7] // U+826F <cjk>
	`諒`: [u8(0x97), 0xC8] // U+8AD2 <cjk>
	`遼`: [u8(0x97), 0xC9] // U+907C <cjk>
	`量`: [u8(0x97), 0xCA] // U+91CF <cjk>
	`陵`: [u8(0x97), 0xCB] // U+9675 <cjk>
	`領`: [u8(0x97), 0xCC] // U+9818 <cjk>
	`力`: [u8(0x97), 0xCD] // U+529B <cjk>
	`緑`: [u8(0x97), 0xCE] // U+7DD1 <cjk>
	`倫`: [u8(0x97), 0xCF] // U+502B <cjk>
	`厘`: [u8(0x97), 0xD0] // U+5398 <cjk>
	`林`: [u8(0x97), 0xD1] // U+6797 <cjk>
	`淋`: [u8(0x97), 0xD2] // U+6DCB <cjk>
	`燐`: [u8(0x97), 0xD3] // U+71D0 <cjk>
	`琳`: [u8(0x97), 0xD4] // U+7433 <cjk>
	`臨`: [u8(0x97), 0xD5] // U+81E8 <cjk>
	`輪`: [u8(0x97), 0xD6] // U+8F2A <cjk>
	`隣`: [u8(0x97), 0xD7] // U+96A3 <cjk>
	`鱗`: [u8(0x97), 0xD8] // U+9C57 <cjk>
	`麟`: [u8(0x97), 0xD9] // U+9E9F <cjk>
	`瑠`: [u8(0x97), 0xDA] // U+7460 <cjk>
	`塁`: [u8(0x97), 0xDB] // U+5841 <cjk>
	`涙`: [u8(0x97), 0xDC] // U+6D99 <cjk>
	`累`: [u8(0x97), 0xDD] // U+7D2F <cjk>
	`類`: [u8(0x97), 0xDE] // U+985E <cjk>
	`令`: [u8(0x97), 0xDF] // U+4EE4 <cjk>
	`伶`: [u8(0x97), 0xE0] // U+4F36 <cjk>
	`例`: [u8(0x97), 0xE1] // U+4F8B <cjk>
	`冷`: [u8(0x97), 0xE2] // U+51B7 <cjk>
	`励`: [u8(0x97), 0xE3] // U+52B1 <cjk>
	`嶺`: [u8(0x97), 0xE4] // U+5DBA <cjk>
	`怜`: [u8(0x97), 0xE5] // U+601C <cjk>
	`玲`: [u8(0x97), 0xE6] // U+73B2 <cjk>
	`礼`: [u8(0x97), 0xE7] // U+793C <cjk>
	`苓`: [u8(0x97), 0xE8] // U+82D3 <cjk>
	`鈴`: [u8(0x97), 0xE9] // U+9234 <cjk>
	`隷`: [u8(0x97), 0xEA] // U+96B7 <cjk>
	`零`: [u8(0x97), 0xEB] // U+96F6 <cjk>
	`霊`: [u8(0x97), 0xEC] // U+970A <cjk>
	`麗`: [u8(0x97), 0xED] // U+9E97 <cjk>
	`齢`: [u8(0x97), 0xEE] // U+9F62 <cjk>
	`暦`: [u8(0x97), 0xEF] // U+66A6 <cjk>
	`歴`: [u8(0x97), 0xF0] // U+6B74 <cjk>
	`列`: [u8(0x97), 0xF1] // U+5217 <cjk>
	`劣`: [u8(0x97), 0xF2] // U+52A3 <cjk>
	`烈`: [u8(0x97), 0xF3] // U+70C8 <cjk>
	`裂`: [u8(0x97), 0xF4] // U+88C2 <cjk>
	`廉`: [u8(0x97), 0xF5] // U+5EC9 <cjk>
	`恋`: [u8(0x97), 0xF6] // U+604B <cjk>
	`憐`: [u8(0x97), 0xF7] // U+6190 <cjk>
	`漣`: [u8(0x97), 0xF8] // U+6F23 <cjk>
	`煉`: [u8(0x97), 0xF9] // U+7149 <cjk>
	`簾`: [u8(0x97), 0xFA] // U+7C3E <cjk>
	`練`: [u8(0x97), 0xFB] // U+7DF4 <cjk>
	`聯`: [u8(0x97), 0xFC] // U+806F <cjk>
	`蓮`: [u8(0x98), 0x40] // U+84EE <cjk>
	`連`: [u8(0x98), 0x41] // U+9023 <cjk>
	`錬`: [u8(0x98), 0x42] // U+932C <cjk>
	`呂`: [u8(0x98), 0x43] // U+5442 <cjk>
	`魯`: [u8(0x98), 0x44] // U+9B6F <cjk>
	`櫓`: [u8(0x98), 0x45] // U+6AD3 <cjk>
	`炉`: [u8(0x98), 0x46] // U+7089 <cjk>
	`賂`: [u8(0x98), 0x47] // U+8CC2 <cjk>
	`路`: [u8(0x98), 0x48] // U+8DEF <cjk>
	`露`: [u8(0x98), 0x49] // U+9732 <cjk>
	`労`: [u8(0x98), 0x4A] // U+52B4 <cjk>
	`婁`: [u8(0x98), 0x4B] // U+5A41 <cjk>
	`廊`: [u8(0x98), 0x4C] // U+5ECA <cjk>
	`弄`: [u8(0x98), 0x4D] // U+5F04 <cjk>
	`朗`: [u8(0x98), 0x4E] // U+6717 <cjk>
	`楼`: [u8(0x98), 0x4F] // U+697C <cjk>
	`榔`: [u8(0x98), 0x50] // U+6994 <cjk>
	`浪`: [u8(0x98), 0x51] // U+6D6A <cjk>
	`漏`: [u8(0x98), 0x52] // U+6F0F <cjk>
	`牢`: [u8(0x98), 0x53] // U+7262 <cjk>
	`狼`: [u8(0x98), 0x54] // U+72FC <cjk>
	`篭`: [u8(0x98), 0x55] // U+7BED <cjk>
	`老`: [u8(0x98), 0x56] // U+8001 <cjk>
	`聾`: [u8(0x98), 0x57] // U+807E <cjk>
	`蝋`: [u8(0x98), 0x58] // U+874B <cjk>
	`郎`: [u8(0x98), 0x59] // U+90CE <cjk>
	`六`: [u8(0x98), 0x5A] // U+516D <cjk>
	`麓`: [u8(0x98), 0x5B] // U+9E93 <cjk>
	`禄`: [u8(0x98), 0x5C] // U+7984 <cjk>
	`肋`: [u8(0x98), 0x5D] // U+808B <cjk>
	`録`: [u8(0x98), 0x5E] // U+9332 <cjk>
	`論`: [u8(0x98), 0x5F] // U+8AD6 <cjk>
	`倭`: [u8(0x98), 0x60] // U+502D <cjk>
	`和`: [u8(0x98), 0x61] // U+548C <cjk>
	`話`: [u8(0x98), 0x62] // U+8A71 <cjk>
	`歪`: [u8(0x98), 0x63] // U+6B6A <cjk>
	`賄`: [u8(0x98), 0x64] // U+8CC4 <cjk>
	`脇`: [u8(0x98), 0x65] // U+8107 <cjk>
	`惑`: [u8(0x98), 0x66] // U+60D1 <cjk>
	`枠`: [u8(0x98), 0x67] // U+67A0 <cjk>
	`鷲`: [u8(0x98), 0x68] // U+9DF2 <cjk>
	`亙`: [u8(0x98), 0x69] // U+4E99 <cjk>
	`亘`: [u8(0x98), 0x6A] // U+4E98 <cjk>
	`鰐`: [u8(0x98), 0x6B] // U+9C10 <cjk>
	`詫`: [u8(0x98), 0x6C] // U+8A6B <cjk>
	`藁`: [u8(0x98), 0x6D] // U+85C1 <cjk>
	`蕨`: [u8(0x98), 0x6E] // U+8568 <cjk>
	`椀`: [u8(0x98), 0x6F] // U+6900 <cjk>
	`湾`: [u8(0x98), 0x70] // U+6E7E <cjk>
	`碗`: [u8(0x98), 0x71] // U+7897 <cjk>
	`腕`: [u8(0x98), 0x72] // U+8155 <cjk>
	`𠮟`: [u8(0x98), 0x73] // U+20B9F <cjk>
	`孁`: [u8(0x98), 0x74] // U+5B41 <cjk>
	`孖`: [u8(0x98), 0x75] // U+5B56 <cjk>
	`孽`: [u8(0x98), 0x76] // U+5B7D <cjk>
	`宓`: [u8(0x98), 0x77] // U+5B93 <cjk>
	`寘`: [u8(0x98), 0x78] // U+5BD8 <cjk>
	`寬`: [u8(0x98), 0x79] // U+5BEC <cjk>
	`尒`: [u8(0x98), 0x7A] // U+5C12 <cjk>
	`尞`: [u8(0x98), 0x7B] // U+5C1E <cjk>
	`尣`: [u8(0x98), 0x7C] // U+5C23 <cjk>
	`尫`: [u8(0x98), 0x7D] // U+5C2B <cjk>
	`㞍`: [u8(0x98), 0x7E] // U+378D <cjk>
	`屢`: [u8(0x98), 0x80] // U+5C62 <cjk>
	`層`: [u8(0x98), 0x81] // U+FA3B CJK COMPATIBILITY IDEOGRAPH-FA3B
	`屮`: [u8(0x98), 0x82] // U+FA3C CJK COMPATIBILITY IDEOGRAPH-FA3C
	`𡚴`: [u8(0x98), 0x83] // U+216B4 <cjk>
	`屺`: [u8(0x98), 0x84] // U+5C7A <cjk>
	`岏`: [u8(0x98), 0x85] // U+5C8F <cjk>
	`岟`: [u8(0x98), 0x86] // U+5C9F <cjk>
	`岣`: [u8(0x98), 0x87] // U+5CA3 <cjk>
	`岪`: [u8(0x98), 0x88] // U+5CAA <cjk>
	`岺`: [u8(0x98), 0x89] // U+5CBA <cjk>
	`峋`: [u8(0x98), 0x8A] // U+5CCB <cjk>
	`峐`: [u8(0x98), 0x8B] // U+5CD0 <cjk>
	`峒`: [u8(0x98), 0x8C] // U+5CD2 <cjk>
	`峴`: [u8(0x98), 0x8D] // U+5CF4 <cjk>
	`𡸴`: [u8(0x98), 0x8E] // U+21E34 <cjk>
	`㟢`: [u8(0x98), 0x8F] // U+37E2 <cjk>
	`崍`: [u8(0x98), 0x90] // U+5D0D <cjk>
	`崧`: [u8(0x98), 0x91] // U+5D27 <cjk>
	`﨑`: [u8(0x98), 0x92] // U+FA11 CJK COMPATIBILITY IDEOGRAPH-FA11
	`嵆`: [u8(0x98), 0x93] // U+5D46 <cjk>
	`嵇`: [u8(0x98), 0x94] // U+5D47 <cjk>
	`嵓`: [u8(0x98), 0x95] // U+5D53 <cjk>
	`嵊`: [u8(0x98), 0x96] // U+5D4A <cjk>
	`嵭`: [u8(0x98), 0x97] // U+5D6D <cjk>
	`嶁`: [u8(0x98), 0x98] // U+5D81 <cjk>
	`嶠`: [u8(0x98), 0x99] // U+5DA0 <cjk>
	`嶤`: [u8(0x98), 0x9A] // U+5DA4 <cjk>
	`嶧`: [u8(0x98), 0x9B] // U+5DA7 <cjk>
	`嶸`: [u8(0x98), 0x9C] // U+5DB8 <cjk>
	`巋`: [u8(0x98), 0x9D] // U+5DCB <cjk>
	`吞`: [u8(0x98), 0x9E] // U+541E <cjk>
	`弌`: [u8(0x98), 0x9F] // U+5F0C <cjk>
	`丐`: [u8(0x98), 0xA0] // U+4E10 <cjk>
	`丕`: [u8(0x98), 0xA1] // U+4E15 <cjk>
	`个`: [u8(0x98), 0xA2] // U+4E2A <cjk>
	`丱`: [u8(0x98), 0xA3] // U+4E31 <cjk>
	`丶`: [u8(0x98), 0xA4] // U+4E36 <cjk>
	`丼`: [u8(0x98), 0xA5] // U+4E3C <cjk>
	`丿`: [u8(0x98), 0xA6] // U+4E3F <cjk>
	`乂`: [u8(0x98), 0xA7] // U+4E42 <cjk>
	`乖`: [u8(0x98), 0xA8] // U+4E56 <cjk>
	`乘`: [u8(0x98), 0xA9] // U+4E58 <cjk>
	`亂`: [u8(0x98), 0xAA] // U+4E82 <cjk>
	`亅`: [u8(0x98), 0xAB] // U+4E85 <cjk>
	`豫`: [u8(0x98), 0xAC] // U+8C6B <cjk>
	`亊`: [u8(0x98), 0xAD] // U+4E8A <cjk>
	`舒`: [u8(0x98), 0xAE] // U+8212 <cjk>
	`弍`: [u8(0x98), 0xAF] // U+5F0D <cjk>
	`于`: [u8(0x98), 0xB0] // U+4E8E <cjk>
	`亞`: [u8(0x98), 0xB1] // U+4E9E <cjk>
	`亟`: [u8(0x98), 0xB2] // U+4E9F <cjk>
	`亠`: [u8(0x98), 0xB3] // U+4EA0 <cjk>
	`亢`: [u8(0x98), 0xB4] // U+4EA2 <cjk>
	`亰`: [u8(0x98), 0xB5] // U+4EB0 <cjk>
	`亳`: [u8(0x98), 0xB6] // U+4EB3 <cjk>
	`亶`: [u8(0x98), 0xB7] // U+4EB6 <cjk>
	`从`: [u8(0x98), 0xB8] // U+4ECE <cjk>
	`仍`: [u8(0x98), 0xB9] // U+4ECD <cjk>
	`仄`: [u8(0x98), 0xBA] // U+4EC4 <cjk>
	`仆`: [u8(0x98), 0xBB] // U+4EC6 <cjk>
	`仂`: [u8(0x98), 0xBC] // U+4EC2 <cjk>
	`仗`: [u8(0x98), 0xBD] // U+4ED7 <cjk>
	`仞`: [u8(0x98), 0xBE] // U+4EDE <cjk>
	`仭`: [u8(0x98), 0xBF] // U+4EED <cjk>
	`仟`: [u8(0x98), 0xC0] // U+4EDF <cjk>
	`价`: [u8(0x98), 0xC1] // U+4EF7 <cjk>
	`伉`: [u8(0x98), 0xC2] // U+4F09 <cjk>
	`佚`: [u8(0x98), 0xC3] // U+4F5A <cjk>
	`估`: [u8(0x98), 0xC4] // U+4F30 <cjk>
	`佛`: [u8(0x98), 0xC5] // U+4F5B <cjk>
	`佝`: [u8(0x98), 0xC6] // U+4F5D <cjk>
	`佗`: [u8(0x98), 0xC7] // U+4F57 <cjk>
	`佇`: [u8(0x98), 0xC8] // U+4F47 <cjk>
	`佶`: [u8(0x98), 0xC9] // U+4F76 <cjk>
	`侈`: [u8(0x98), 0xCA] // U+4F88 <cjk>
	`侏`: [u8(0x98), 0xCB] // U+4F8F <cjk>
	`侘`: [u8(0x98), 0xCC] // U+4F98 <cjk>
	`佻`: [u8(0x98), 0xCD] // U+4F7B <cjk>
	`佩`: [u8(0x98), 0xCE] // U+4F69 <cjk>
	`佰`: [u8(0x98), 0xCF] // U+4F70 <cjk>
	`侑`: [u8(0x98), 0xD0] // U+4F91 <cjk>
	`佯`: [u8(0x98), 0xD1] // U+4F6F <cjk>
	`來`: [u8(0x98), 0xD2] // U+4F86 <cjk>
	`侖`: [u8(0x98), 0xD3] // U+4F96 <cjk>
	`儘`: [u8(0x98), 0xD4] // U+5118 <cjk>
	`俔`: [u8(0x98), 0xD5] // U+4FD4 <cjk>
	`俟`: [u8(0x98), 0xD6] // U+4FDF <cjk>
	`俎`: [u8(0x98), 0xD7] // U+4FCE <cjk>
	`俘`: [u8(0x98), 0xD8] // U+4FD8 <cjk>
	`俛`: [u8(0x98), 0xD9] // U+4FDB <cjk>
	`俑`: [u8(0x98), 0xDA] // U+4FD1 <cjk>
	`俚`: [u8(0x98), 0xDB] // U+4FDA <cjk>
	`俐`: [u8(0x98), 0xDC] // U+4FD0 <cjk>
	`俤`: [u8(0x98), 0xDD] // U+4FE4 <cjk>
	`俥`: [u8(0x98), 0xDE] // U+4FE5 <cjk>
	`倚`: [u8(0x98), 0xDF] // U+501A <cjk>
	`倨`: [u8(0x98), 0xE0] // U+5028 <cjk>
	`倔`: [u8(0x98), 0xE1] // U+5014 <cjk>
	`倪`: [u8(0x98), 0xE2] // U+502A <cjk>
	`倥`: [u8(0x98), 0xE3] // U+5025 <cjk>
	`倅`: [u8(0x98), 0xE4] // U+5005 <cjk>
	`伜`: [u8(0x98), 0xE5] // U+4F1C <cjk>
	`俶`: [u8(0x98), 0xE6] // U+4FF6 <cjk>
	`倡`: [u8(0x98), 0xE7] // U+5021 <cjk>
	`倩`: [u8(0x98), 0xE8] // U+5029 <cjk>
	`倬`: [u8(0x98), 0xE9] // U+502C <cjk>
	`俾`: [u8(0x98), 0xEA] // U+4FFE <cjk>
	`俯`: [u8(0x98), 0xEB] // U+4FEF <cjk>
	`們`: [u8(0x98), 0xEC] // U+5011 <cjk>
	`倆`: [u8(0x98), 0xED] // U+5006 <cjk>
	`偃`: [u8(0x98), 0xEE] // U+5043 <cjk>
	`假`: [u8(0x98), 0xEF] // U+5047 <cjk>
	`會`: [u8(0x98), 0xF0] // U+6703 <cjk>
	`偕`: [u8(0x98), 0xF1] // U+5055 <cjk>
	`偐`: [u8(0x98), 0xF2] // U+5050 <cjk>
	`偈`: [u8(0x98), 0xF3] // U+5048 <cjk>
	`做`: [u8(0x98), 0xF4] // U+505A <cjk>
	`偖`: [u8(0x98), 0xF5] // U+5056 <cjk>
	`偬`: [u8(0x98), 0xF6] // U+506C <cjk>
	`偸`: [u8(0x98), 0xF7] // U+5078 <cjk>
	`傀`: [u8(0x98), 0xF8] // U+5080 <cjk>
	`傚`: [u8(0x98), 0xF9] // U+509A <cjk>
	`傅`: [u8(0x98), 0xFA] // U+5085 <cjk>
	`傴`: [u8(0x98), 0xFB] // U+50B4 <cjk>
	`傲`: [u8(0x98), 0xFC] // U+50B2 <cjk>
	`僉`: [u8(0x99), 0x40] // U+50C9 <cjk>
	`僊`: [u8(0x99), 0x41] // U+50CA <cjk>
	`傳`: [u8(0x99), 0x42] // U+50B3 <cjk>
	`僂`: [u8(0x99), 0x43] // U+50C2 <cjk>
	`僖`: [u8(0x99), 0x44] // U+50D6 <cjk>
	`僞`: [u8(0x99), 0x45] // U+50DE <cjk>
	`僥`: [u8(0x99), 0x46] // U+50E5 <cjk>
	`僭`: [u8(0x99), 0x47] // U+50ED <cjk>
	`僣`: [u8(0x99), 0x48] // U+50E3 <cjk>
	`僮`: [u8(0x99), 0x49] // U+50EE <cjk>
	`價`: [u8(0x99), 0x4A] // U+50F9 <cjk>
	`僵`: [u8(0x99), 0x4B] // U+50F5 <cjk>
	`儉`: [u8(0x99), 0x4C] // U+5109 <cjk>
	`儁`: [u8(0x99), 0x4D] // U+5101 <cjk>
	`儂`: [u8(0x99), 0x4E] // U+5102 <cjk>
	`儖`: [u8(0x99), 0x4F] // U+5116 <cjk>
	`儕`: [u8(0x99), 0x50] // U+5115 <cjk>
	`儔`: [u8(0x99), 0x51] // U+5114 <cjk>
	`儚`: [u8(0x99), 0x52] // U+511A <cjk>
	`儡`: [u8(0x99), 0x53] // U+5121 <cjk>
	`儺`: [u8(0x99), 0x54] // U+513A <cjk>
	`儷`: [u8(0x99), 0x55] // U+5137 <cjk>
	`儼`: [u8(0x99), 0x56] // U+513C <cjk>
	`儻`: [u8(0x99), 0x57] // U+513B <cjk>
	`儿`: [u8(0x99), 0x58] // U+513F <cjk>
	`兀`: [u8(0x99), 0x59] // U+5140 <cjk>
	`兒`: [u8(0x99), 0x5A] // U+5152 <cjk>
	`兌`: [u8(0x99), 0x5B] // U+514C <cjk>
	`兔`: [u8(0x99), 0x5C] // U+5154 <cjk>
	`兢`: [u8(0x99), 0x5D] // U+5162 <cjk>
	`竸`: [u8(0x99), 0x5E] // U+7AF8 <cjk>
	`兩`: [u8(0x99), 0x5F] // U+5169 <cjk>
	`兪`: [u8(0x99), 0x60] // U+516A <cjk>
	`兮`: [u8(0x99), 0x61] // U+516E <cjk>
	`冀`: [u8(0x99), 0x62] // U+5180 <cjk>
	`冂`: [u8(0x99), 0x63] // U+5182 <cjk>
	`囘`: [u8(0x99), 0x64] // U+56D8 <cjk>
	`册`: [u8(0x99), 0x65] // U+518C <cjk>
	`冉`: [u8(0x99), 0x66] // U+5189 <cjk>
	`冏`: [u8(0x99), 0x67] // U+518F <cjk>
	`冑`: [u8(0x99), 0x68] // U+5191 <cjk>
	`冓`: [u8(0x99), 0x69] // U+5193 <cjk>
	`冕`: [u8(0x99), 0x6A] // U+5195 <cjk>
	`冖`: [u8(0x99), 0x6B] // U+5196 <cjk>
	`冤`: [u8(0x99), 0x6C] // U+51A4 <cjk>
	`冦`: [u8(0x99), 0x6D] // U+51A6 <cjk>
	`冢`: [u8(0x99), 0x6E] // U+51A2 <cjk>
	`冩`: [u8(0x99), 0x6F] // U+51A9 <cjk>
	`冪`: [u8(0x99), 0x70] // U+51AA <cjk>
	`冫`: [u8(0x99), 0x71] // U+51AB <cjk>
	`决`: [u8(0x99), 0x72] // U+51B3 <cjk>
	`冱`: [u8(0x99), 0x73] // U+51B1 <cjk>
	`冲`: [u8(0x99), 0x74] // U+51B2 <cjk>
	`冰`: [u8(0x99), 0x75] // U+51B0 <cjk>
	`况`: [u8(0x99), 0x76] // U+51B5 <cjk>
	`冽`: [u8(0x99), 0x77] // U+51BD <cjk>
	`凅`: [u8(0x99), 0x78] // U+51C5 <cjk>
	`凉`: [u8(0x99), 0x79] // U+51C9 <cjk>
	`凛`: [u8(0x99), 0x7A] // U+51DB <cjk>
	`几`: [u8(0x99), 0x7B] // U+51E0 <cjk>
	`處`: [u8(0x99), 0x7C] // U+8655 <cjk>
	`凩`: [u8(0x99), 0x7D] // U+51E9 <cjk>
	`凭`: [u8(0x99), 0x7E] // U+51ED <cjk>
	`凰`: [u8(0x99), 0x80] // U+51F0 <cjk>
	`凵`: [u8(0x99), 0x81] // U+51F5 <cjk>
	`凾`: [u8(0x99), 0x82] // U+51FE <cjk>
	`刄`: [u8(0x99), 0x83] // U+5204 <cjk>
	`刋`: [u8(0x99), 0x84] // U+520B <cjk>
	`刔`: [u8(0x99), 0x85] // U+5214 <cjk>
	`刎`: [u8(0x99), 0x86] // U+520E <cjk>
	`刧`: [u8(0x99), 0x87] // U+5227 <cjk>
	`刪`: [u8(0x99), 0x88] // U+522A <cjk>
	`刮`: [u8(0x99), 0x89] // U+522E <cjk>
	`刳`: [u8(0x99), 0x8A] // U+5233 <cjk>
	`刹`: [u8(0x99), 0x8B] // U+5239 <cjk>
	`剏`: [u8(0x99), 0x8C] // U+524F <cjk>
	`剄`: [u8(0x99), 0x8D] // U+5244 <cjk>
	`剋`: [u8(0x99), 0x8E] // U+524B <cjk>
	`剌`: [u8(0x99), 0x8F] // U+524C <cjk>
	`剞`: [u8(0x99), 0x90] // U+525E <cjk>
	`剔`: [u8(0x99), 0x91] // U+5254 <cjk>
	`剪`: [u8(0x99), 0x92] // U+526A <cjk>
	`剴`: [u8(0x99), 0x93] // U+5274 <cjk>
	`剩`: [u8(0x99), 0x94] // U+5269 <cjk>
	`剳`: [u8(0x99), 0x95] // U+5273 <cjk>
	`剿`: [u8(0x99), 0x96] // U+527F <cjk>
	`剽`: [u8(0x99), 0x97] // U+527D <cjk>
	`劍`: [u8(0x99), 0x98] // U+528D <cjk>
	`劔`: [u8(0x99), 0x99] // U+5294 <cjk>
	`劒`: [u8(0x99), 0x9A] // U+5292 <cjk>
	`剱`: [u8(0x99), 0x9B] // U+5271 <cjk>
	`劈`: [u8(0x99), 0x9C] // U+5288 <cjk>
	`劑`: [u8(0x99), 0x9D] // U+5291 <cjk>
	`辨`: [u8(0x99), 0x9E] // U+8FA8 <cjk>
	`辧`: [u8(0x99), 0x9F] // U+8FA7 <cjk>
	`劬`: [u8(0x99), 0xA0] // U+52AC <cjk>
	`劭`: [u8(0x99), 0xA1] // U+52AD <cjk>
	`劼`: [u8(0x99), 0xA2] // U+52BC <cjk>
	`劵`: [u8(0x99), 0xA3] // U+52B5 <cjk>
	`勁`: [u8(0x99), 0xA4] // U+52C1 <cjk>
	`勍`: [u8(0x99), 0xA5] // U+52CD <cjk>
	`勗`: [u8(0x99), 0xA6] // U+52D7 <cjk>
	`勞`: [u8(0x99), 0xA7] // U+52DE <cjk>
	`勣`: [u8(0x99), 0xA8] // U+52E3 <cjk>
	`勦`: [u8(0x99), 0xA9] // U+52E6 <cjk>
	`飭`: [u8(0x99), 0xAA] // U+98ED <cjk>
	`勠`: [u8(0x99), 0xAB] // U+52E0 <cjk>
	`勳`: [u8(0x99), 0xAC] // U+52F3 <cjk>
	`勵`: [u8(0x99), 0xAD] // U+52F5 <cjk>
	`勸`: [u8(0x99), 0xAE] // U+52F8 <cjk>
	`勹`: [u8(0x99), 0xAF] // U+52F9 <cjk>
	`匆`: [u8(0x99), 0xB0] // U+5306 <cjk>
	`匈`: [u8(0x99), 0xB1] // U+5308 <cjk>
	`甸`: [u8(0x99), 0xB2] // U+7538 <cjk>
	`匍`: [u8(0x99), 0xB3] // U+530D <cjk>
	`匐`: [u8(0x99), 0xB4] // U+5310 <cjk>
	`匏`: [u8(0x99), 0xB5] // U+530F <cjk>
	`匕`: [u8(0x99), 0xB6] // U+5315 <cjk>
	`匚`: [u8(0x99), 0xB7] // U+531A <cjk>
	`匣`: [u8(0x99), 0xB8] // U+5323 <cjk>
	`匯`: [u8(0x99), 0xB9] // U+532F <cjk>
	`匱`: [u8(0x99), 0xBA] // U+5331 <cjk>
	`匳`: [u8(0x99), 0xBB] // U+5333 <cjk>
	`匸`: [u8(0x99), 0xBC] // U+5338 <cjk>
	`區`: [u8(0x99), 0xBD] // U+5340 <cjk>
	`卆`: [u8(0x99), 0xBE] // U+5346 <cjk>
	`卅`: [u8(0x99), 0xBF] // U+5345 <cjk>
	`丗`: [u8(0x99), 0xC0] // U+4E17 <cjk>
	`卉`: [u8(0x99), 0xC1] // U+5349 <cjk>
	`卍`: [u8(0x99), 0xC2] // U+534D <cjk>
	`凖`: [u8(0x99), 0xC3] // U+51D6 <cjk>
	`卞`: [u8(0x99), 0xC4] // U+535E <cjk>
	`卩`: [u8(0x99), 0xC5] // U+5369 <cjk>
	`卮`: [u8(0x99), 0xC6] // U+536E <cjk>
	`夘`: [u8(0x99), 0xC7] // U+5918 <cjk>
	`卻`: [u8(0x99), 0xC8] // U+537B <cjk>
	`卷`: [u8(0x99), 0xC9] // U+5377 <cjk>
	`厂`: [u8(0x99), 0xCA] // U+5382 <cjk>
	`厖`: [u8(0x99), 0xCB] // U+5396 <cjk>
	`厠`: [u8(0x99), 0xCC] // U+53A0 <cjk>
	`厦`: [u8(0x99), 0xCD] // U+53A6 <cjk>
	`厥`: [u8(0x99), 0xCE] // U+53A5 <cjk>
	`厮`: [u8(0x99), 0xCF] // U+53AE <cjk>
	`厰`: [u8(0x99), 0xD0] // U+53B0 <cjk>
	`厶`: [u8(0x99), 0xD1] // U+53B6 <cjk>
	`參`: [u8(0x99), 0xD2] // U+53C3 <cjk>
	`簒`: [u8(0x99), 0xD3] // U+7C12 <cjk>
	`雙`: [u8(0x99), 0xD4] // U+96D9 <cjk>
	`叟`: [u8(0x99), 0xD5] // U+53DF <cjk>
	`曼`: [u8(0x99), 0xD6] // U+66FC <cjk>
	`燮`: [u8(0x99), 0xD7] // U+71EE <cjk>
	`叮`: [u8(0x99), 0xD8] // U+53EE <cjk>
	`叨`: [u8(0x99), 0xD9] // U+53E8 <cjk>
	`叭`: [u8(0x99), 0xDA] // U+53ED <cjk>
	`叺`: [u8(0x99), 0xDB] // U+53FA <cjk>
	`吁`: [u8(0x99), 0xDC] // U+5401 <cjk>
	`吽`: [u8(0x99), 0xDD] // U+543D <cjk>
	`呀`: [u8(0x99), 0xDE] // U+5440 <cjk>
	`听`: [u8(0x99), 0xDF] // U+542C <cjk>
	`吭`: [u8(0x99), 0xE0] // U+542D <cjk>
	`吼`: [u8(0x99), 0xE1] // U+543C <cjk>
	`吮`: [u8(0x99), 0xE2] // U+542E <cjk>
	`吶`: [u8(0x99), 0xE3] // U+5436 <cjk>
	`吩`: [u8(0x99), 0xE4] // U+5429 <cjk>
	`吝`: [u8(0x99), 0xE5] // U+541D <cjk>
	`呎`: [u8(0x99), 0xE6] // U+544E <cjk>
	`咏`: [u8(0x99), 0xE7] // U+548F <cjk>
	`呵`: [u8(0x99), 0xE8] // U+5475 <cjk>
	`咎`: [u8(0x99), 0xE9] // U+548E <cjk>
	`呟`: [u8(0x99), 0xEA] // U+545F <cjk>
	`呱`: [u8(0x99), 0xEB] // U+5471 <cjk>
	`呷`: [u8(0x99), 0xEC] // U+5477 <cjk>
	`呰`: [u8(0x99), 0xED] // U+5470 <cjk>
	`咒`: [u8(0x99), 0xEE] // U+5492 <cjk>
	`呻`: [u8(0x99), 0xEF] // U+547B <cjk>
	`咀`: [u8(0x99), 0xF0] // U+5480 <cjk>
	`呶`: [u8(0x99), 0xF1] // U+5476 <cjk>
	`咄`: [u8(0x99), 0xF2] // U+5484 <cjk>
	`咐`: [u8(0x99), 0xF3] // U+5490 <cjk>
	`咆`: [u8(0x99), 0xF4] // U+5486 <cjk>
	`哇`: [u8(0x99), 0xF5] // U+54C7 <cjk>
	`咢`: [u8(0x99), 0xF6] // U+54A2 <cjk>
	`咸`: [u8(0x99), 0xF7] // U+54B8 <cjk>
	`咥`: [u8(0x99), 0xF8] // U+54A5 <cjk>
	`咬`: [u8(0x99), 0xF9] // U+54AC <cjk>
	`哄`: [u8(0x99), 0xFA] // U+54C4 <cjk>
	`哈`: [u8(0x99), 0xFB] // U+54C8 <cjk>
	`咨`: [u8(0x99), 0xFC] // U+54A8 <cjk>
	`咫`: [u8(0x9A), 0x40] // U+54AB <cjk>
	`哂`: [u8(0x9A), 0x41] // U+54C2 <cjk>
	`咤`: [u8(0x9A), 0x42] // U+54A4 <cjk>
	`咾`: [u8(0x9A), 0x43] // U+54BE <cjk>
	`咼`: [u8(0x9A), 0x44] // U+54BC <cjk>
	`哘`: [u8(0x9A), 0x45] // U+54D8 <cjk>
	`哥`: [u8(0x9A), 0x46] // U+54E5 <cjk>
	`哦`: [u8(0x9A), 0x47] // U+54E6 <cjk>
	`唏`: [u8(0x9A), 0x48] // U+550F <cjk>
	`唔`: [u8(0x9A), 0x49] // U+5514 <cjk>
	`哽`: [u8(0x9A), 0x4A] // U+54FD <cjk>
	`哮`: [u8(0x9A), 0x4B] // U+54EE <cjk>
	`哭`: [u8(0x9A), 0x4C] // U+54ED <cjk>
	`哺`: [u8(0x9A), 0x4D] // U+54FA <cjk>
	`哢`: [u8(0x9A), 0x4E] // U+54E2 <cjk>
	`唹`: [u8(0x9A), 0x4F] // U+5539 <cjk>
	`啀`: [u8(0x9A), 0x50] // U+5540 <cjk>
	`啣`: [u8(0x9A), 0x51] // U+5563 <cjk>
	`啌`: [u8(0x9A), 0x52] // U+554C <cjk>
	`售`: [u8(0x9A), 0x53] // U+552E <cjk>
	`啜`: [u8(0x9A), 0x54] // U+555C <cjk>
	`啅`: [u8(0x9A), 0x55] // U+5545 <cjk>
	`啖`: [u8(0x9A), 0x56] // U+5556 <cjk>
	`啗`: [u8(0x9A), 0x57] // U+5557 <cjk>
	`唸`: [u8(0x9A), 0x58] // U+5538 <cjk>
	`唳`: [u8(0x9A), 0x59] // U+5533 <cjk>
	`啝`: [u8(0x9A), 0x5A] // U+555D <cjk>
	`喙`: [u8(0x9A), 0x5B] // U+5599 <cjk>
	`喀`: [u8(0x9A), 0x5C] // U+5580 <cjk>
	`咯`: [u8(0x9A), 0x5D] // U+54AF <cjk>
	`喊`: [u8(0x9A), 0x5E] // U+558A <cjk>
	`喟`: [u8(0x9A), 0x5F] // U+559F <cjk>
	`啻`: [u8(0x9A), 0x60] // U+557B <cjk>
	`啾`: [u8(0x9A), 0x61] // U+557E <cjk>
	`喘`: [u8(0x9A), 0x62] // U+5598 <cjk>
	`喞`: [u8(0x9A), 0x63] // U+559E <cjk>
	`單`: [u8(0x9A), 0x64] // U+55AE <cjk>
	`啼`: [u8(0x9A), 0x65] // U+557C <cjk>
	`喃`: [u8(0x9A), 0x66] // U+5583 <cjk>
	`喩`: [u8(0x9A), 0x67] // U+55A9 <cjk>
	`喇`: [u8(0x9A), 0x68] // U+5587 <cjk>
	`喨`: [u8(0x9A), 0x69] // U+55A8 <cjk>
	`嗚`: [u8(0x9A), 0x6A] // U+55DA <cjk>
	`嗅`: [u8(0x9A), 0x6B] // U+55C5 <cjk>
	`嗟`: [u8(0x9A), 0x6C] // U+55DF <cjk>
	`嗄`: [u8(0x9A), 0x6D] // U+55C4 <cjk>
	`嗜`: [u8(0x9A), 0x6E] // U+55DC <cjk>
	`嗤`: [u8(0x9A), 0x6F] // U+55E4 <cjk>
	`嗔`: [u8(0x9A), 0x70] // U+55D4 <cjk>
	`嘔`: [u8(0x9A), 0x71] // U+5614 <cjk>
	`嗷`: [u8(0x9A), 0x72] // U+55F7 <cjk>
	`嘖`: [u8(0x9A), 0x73] // U+5616 <cjk>
	`嗾`: [u8(0x9A), 0x74] // U+55FE <cjk>
	`嗽`: [u8(0x9A), 0x75] // U+55FD <cjk>
	`嘛`: [u8(0x9A), 0x76] // U+561B <cjk>
	`嗹`: [u8(0x9A), 0x77] // U+55F9 <cjk>
	`噎`: [u8(0x9A), 0x78] // U+564E <cjk>
	`噐`: [u8(0x9A), 0x79] // U+5650 <cjk>
	`營`: [u8(0x9A), 0x7A] // U+71DF <cjk>
	`嘴`: [u8(0x9A), 0x7B] // U+5634 <cjk>
	`嘶`: [u8(0x9A), 0x7C] // U+5636 <cjk>
	`嘲`: [u8(0x9A), 0x7D] // U+5632 <cjk>
	`嘸`: [u8(0x9A), 0x7E] // U+5638 <cjk>
	`噫`: [u8(0x9A), 0x80] // U+566B <cjk>
	`噤`: [u8(0x9A), 0x81] // U+5664 <cjk>
	`嘯`: [u8(0x9A), 0x82] // U+562F <cjk>
	`噬`: [u8(0x9A), 0x83] // U+566C <cjk>
	`噪`: [u8(0x9A), 0x84] // U+566A <cjk>
	`嚆`: [u8(0x9A), 0x85] // U+5686 <cjk>
	`嚀`: [u8(0x9A), 0x86] // U+5680 <cjk>
	`嚊`: [u8(0x9A), 0x87] // U+568A <cjk>
	`嚠`: [u8(0x9A), 0x88] // U+56A0 <cjk>
	`嚔`: [u8(0x9A), 0x89] // U+5694 <cjk>
	`嚏`: [u8(0x9A), 0x8A] // U+568F <cjk>
	`嚥`: [u8(0x9A), 0x8B] // U+56A5 <cjk>
	`嚮`: [u8(0x9A), 0x8C] // U+56AE <cjk>
	`嚶`: [u8(0x9A), 0x8D] // U+56B6 <cjk>
	`嚴`: [u8(0x9A), 0x8E] // U+56B4 <cjk>
	`囂`: [u8(0x9A), 0x8F] // U+56C2 <cjk>
	`嚼`: [u8(0x9A), 0x90] // U+56BC <cjk>
	`囁`: [u8(0x9A), 0x91] // U+56C1 <cjk>
	`囃`: [u8(0x9A), 0x92] // U+56C3 <cjk>
	`囀`: [u8(0x9A), 0x93] // U+56C0 <cjk>
	`囈`: [u8(0x9A), 0x94] // U+56C8 <cjk>
	`囎`: [u8(0x9A), 0x95] // U+56CE <cjk>
	`囑`: [u8(0x9A), 0x96] // U+56D1 <cjk>
	`囓`: [u8(0x9A), 0x97] // U+56D3 <cjk>
	`囗`: [u8(0x9A), 0x98] // U+56D7 <cjk>
	`囮`: [u8(0x9A), 0x99] // U+56EE <cjk>
	`囹`: [u8(0x9A), 0x9A] // U+56F9 <cjk>
	`圀`: [u8(0x9A), 0x9B] // U+5700 <cjk>
	`囿`: [u8(0x9A), 0x9C] // U+56FF <cjk>
	`圄`: [u8(0x9A), 0x9D] // U+5704 <cjk>
	`圉`: [u8(0x9A), 0x9E] // U+5709 <cjk>
	`圈`: [u8(0x9A), 0x9F] // U+5708 <cjk>
	`國`: [u8(0x9A), 0xA0] // U+570B <cjk>
	`圍`: [u8(0x9A), 0xA1] // U+570D <cjk>
	`圓`: [u8(0x9A), 0xA2] // U+5713 <cjk>
	`團`: [u8(0x9A), 0xA3] // U+5718 <cjk>
	`圖`: [u8(0x9A), 0xA4] // U+5716 <cjk>
	`嗇`: [u8(0x9A), 0xA5] // U+55C7 <cjk>
	`圜`: [u8(0x9A), 0xA6] // U+571C <cjk>
	`圦`: [u8(0x9A), 0xA7] // U+5726 <cjk>
	`圷`: [u8(0x9A), 0xA8] // U+5737 <cjk>
	`圸`: [u8(0x9A), 0xA9] // U+5738 <cjk>
	`坎`: [u8(0x9A), 0xAA] // U+574E <cjk>
	`圻`: [u8(0x9A), 0xAB] // U+573B <cjk>
	`址`: [u8(0x9A), 0xAC] // U+5740 <cjk>
	`坏`: [u8(0x9A), 0xAD] // U+574F <cjk>
	`坩`: [u8(0x9A), 0xAE] // U+5769 <cjk>
	`埀`: [u8(0x9A), 0xAF] // U+57C0 <cjk>
	`垈`: [u8(0x9A), 0xB0] // U+5788 <cjk>
	`坡`: [u8(0x9A), 0xB1] // U+5761 <cjk>
	`坿`: [u8(0x9A), 0xB2] // U+577F <cjk>
	`垉`: [u8(0x9A), 0xB3] // U+5789 <cjk>
	`垓`: [u8(0x9A), 0xB4] // U+5793 <cjk>
	`垠`: [u8(0x9A), 0xB5] // U+57A0 <cjk>
	`垳`: [u8(0x9A), 0xB6] // U+57B3 <cjk>
	`垤`: [u8(0x9A), 0xB7] // U+57A4 <cjk>
	`垪`: [u8(0x9A), 0xB8] // U+57AA <cjk>
	`垰`: [u8(0x9A), 0xB9] // U+57B0 <cjk>
	`埃`: [u8(0x9A), 0xBA] // U+57C3 <cjk>
	`埆`: [u8(0x9A), 0xBB] // U+57C6 <cjk>
	`埔`: [u8(0x9A), 0xBC] // U+57D4 <cjk>
	`埒`: [u8(0x9A), 0xBD] // U+57D2 <cjk>
	`埓`: [u8(0x9A), 0xBE] // U+57D3 <cjk>
	`堊`: [u8(0x9A), 0xBF] // U+580A <cjk>
	`埖`: [u8(0x9A), 0xC0] // U+57D6 <cjk>
	`埣`: [u8(0x9A), 0xC1] // U+57E3 <cjk>
	`堋`: [u8(0x9A), 0xC2] // U+580B <cjk>
	`堙`: [u8(0x9A), 0xC3] // U+5819 <cjk>
	`堝`: [u8(0x9A), 0xC4] // U+581D <cjk>
	`塲`: [u8(0x9A), 0xC5] // U+5872 <cjk>
	`堡`: [u8(0x9A), 0xC6] // U+5821 <cjk>
	`塢`: [u8(0x9A), 0xC7] // U+5862 <cjk>
	`塋`: [u8(0x9A), 0xC8] // U+584B <cjk>
	`塰`: [u8(0x9A), 0xC9] // U+5870 <cjk>
	`毀`: [u8(0x9A), 0xCA] // U+6BC0 <cjk>
	`塒`: [u8(0x9A), 0xCB] // U+5852 <cjk>
	`堽`: [u8(0x9A), 0xCC] // U+583D <cjk>
	`塹`: [u8(0x9A), 0xCD] // U+5879 <cjk>
	`墅`: [u8(0x9A), 0xCE] // U+5885 <cjk>
	`墹`: [u8(0x9A), 0xCF] // U+58B9 <cjk>
	`墟`: [u8(0x9A), 0xD0] // U+589F <cjk>
	`墫`: [u8(0x9A), 0xD1] // U+58AB <cjk>
	`墺`: [u8(0x9A), 0xD2] // U+58BA <cjk>
	`壞`: [u8(0x9A), 0xD3] // U+58DE <cjk>
	`墻`: [u8(0x9A), 0xD4] // U+58BB <cjk>
	`墸`: [u8(0x9A), 0xD5] // U+58B8 <cjk>
	`墮`: [u8(0x9A), 0xD6] // U+58AE <cjk>
	`壅`: [u8(0x9A), 0xD7] // U+58C5 <cjk>
	`壓`: [u8(0x9A), 0xD8] // U+58D3 <cjk>
	`壑`: [u8(0x9A), 0xD9] // U+58D1 <cjk>
	`壗`: [u8(0x9A), 0xDA] // U+58D7 <cjk>
	`壙`: [u8(0x9A), 0xDB] // U+58D9 <cjk>
	`壘`: [u8(0x9A), 0xDC] // U+58D8 <cjk>
	`壥`: [u8(0x9A), 0xDD] // U+58E5 <cjk>
	`壜`: [u8(0x9A), 0xDE] // U+58DC <cjk>
	`壤`: [u8(0x9A), 0xDF] // U+58E4 <cjk>
	`壟`: [u8(0x9A), 0xE0] // U+58DF <cjk>
	`壯`: [u8(0x9A), 0xE1] // U+58EF <cjk>
	`壺`: [u8(0x9A), 0xE2] // U+58FA <cjk>
	`壹`: [u8(0x9A), 0xE3] // U+58F9 <cjk>
	`壻`: [u8(0x9A), 0xE4] // U+58FB <cjk>
	`壼`: [u8(0x9A), 0xE5] // U+58FC <cjk>
	`壽`: [u8(0x9A), 0xE6] // U+58FD <cjk>
	`夂`: [u8(0x9A), 0xE7] // U+5902 <cjk>
	`夊`: [u8(0x9A), 0xE8] // U+590A <cjk>
	`夐`: [u8(0x9A), 0xE9] // U+5910 <cjk>
	`夛`: [u8(0x9A), 0xEA] // U+591B <cjk>
	`梦`: [u8(0x9A), 0xEB] // U+68A6 <cjk>
	`夥`: [u8(0x9A), 0xEC] // U+5925 <cjk>
	`夬`: [u8(0x9A), 0xED] // U+592C <cjk>
	`夭`: [u8(0x9A), 0xEE] // U+592D <cjk>
	`夲`: [u8(0x9A), 0xEF] // U+5932 <cjk>
	`夸`: [u8(0x9A), 0xF0] // U+5938 <cjk>
	`夾`: [u8(0x9A), 0xF1] // U+593E <cjk>
	`竒`: [u8(0x9A), 0xF2] // U+7AD2 <cjk>
	`奕`: [u8(0x9A), 0xF3] // U+5955 <cjk>
	`奐`: [u8(0x9A), 0xF4] // U+5950 <cjk>
	`奎`: [u8(0x9A), 0xF5] // U+594E <cjk>
	`奚`: [u8(0x9A), 0xF6] // U+595A <cjk>
	`奘`: [u8(0x9A), 0xF7] // U+5958 <cjk>
	`奢`: [u8(0x9A), 0xF8] // U+5962 <cjk>
	`奠`: [u8(0x9A), 0xF9] // U+5960 <cjk>
	`奧`: [u8(0x9A), 0xFA] // U+5967 <cjk>
	`奬`: [u8(0x9A), 0xFB] // U+596C <cjk>
	`奩`: [u8(0x9A), 0xFC] // U+5969 <cjk>
	`奸`: [u8(0x9B), 0x40] // U+5978 <cjk>
	`妁`: [u8(0x9B), 0x41] // U+5981 <cjk>
	`妝`: [u8(0x9B), 0x42] // U+599D <cjk>
	`佞`: [u8(0x9B), 0x43] // U+4F5E <cjk>
	`侫`: [u8(0x9B), 0x44] // U+4FAB <cjk>
	`妣`: [u8(0x9B), 0x45] // U+59A3 <cjk>
	`妲`: [u8(0x9B), 0x46] // U+59B2 <cjk>
	`姆`: [u8(0x9B), 0x47] // U+59C6 <cjk>
	`姨`: [u8(0x9B), 0x48] // U+59E8 <cjk>
	`姜`: [u8(0x9B), 0x49] // U+59DC <cjk>
	`妍`: [u8(0x9B), 0x4A] // U+598D <cjk>
	`姙`: [u8(0x9B), 0x4B] // U+59D9 <cjk>
	`姚`: [u8(0x9B), 0x4C] // U+59DA <cjk>
	`娥`: [u8(0x9B), 0x4D] // U+5A25 <cjk>
	`娟`: [u8(0x9B), 0x4E] // U+5A1F <cjk>
	`娑`: [u8(0x9B), 0x4F] // U+5A11 <cjk>
	`娜`: [u8(0x9B), 0x50] // U+5A1C <cjk>
	`娉`: [u8(0x9B), 0x51] // U+5A09 <cjk>
	`娚`: [u8(0x9B), 0x52] // U+5A1A <cjk>
	`婀`: [u8(0x9B), 0x53] // U+5A40 <cjk>
	`婬`: [u8(0x9B), 0x54] // U+5A6C <cjk>
	`婉`: [u8(0x9B), 0x55] // U+5A49 <cjk>
	`娵`: [u8(0x9B), 0x56] // U+5A35 <cjk>
	`娶`: [u8(0x9B), 0x57] // U+5A36 <cjk>
	`婢`: [u8(0x9B), 0x58] // U+5A62 <cjk>
	`婪`: [u8(0x9B), 0x59] // U+5A6A <cjk>
	`媚`: [u8(0x9B), 0x5A] // U+5A9A <cjk>
	`媼`: [u8(0x9B), 0x5B] // U+5ABC <cjk>
	`媾`: [u8(0x9B), 0x5C] // U+5ABE <cjk>
	`嫋`: [u8(0x9B), 0x5D] // U+5ACB <cjk>
	`嫂`: [u8(0x9B), 0x5E] // U+5AC2 <cjk>
	`媽`: [u8(0x9B), 0x5F] // U+5ABD <cjk>
	`嫣`: [u8(0x9B), 0x60] // U+5AE3 <cjk>
	`嫗`: [u8(0x9B), 0x61] // U+5AD7 <cjk>
	`嫦`: [u8(0x9B), 0x62] // U+5AE6 <cjk>
	`嫩`: [u8(0x9B), 0x63] // U+5AE9 <cjk>
	`嫖`: [u8(0x9B), 0x64] // U+5AD6 <cjk>
	`嫺`: [u8(0x9B), 0x65] // U+5AFA <cjk>
	`嫻`: [u8(0x9B), 0x66] // U+5AFB <cjk>
	`嬌`: [u8(0x9B), 0x67] // U+5B0C <cjk>
	`嬋`: [u8(0x9B), 0x68] // U+5B0B <cjk>
	`嬖`: [u8(0x9B), 0x69] // U+5B16 <cjk>
	`嬲`: [u8(0x9B), 0x6A] // U+5B32 <cjk>
	`嫐`: [u8(0x9B), 0x6B] // U+5AD0 <cjk>
	`嬪`: [u8(0x9B), 0x6C] // U+5B2A <cjk>
	`嬶`: [u8(0x9B), 0x6D] // U+5B36 <cjk>
	`嬾`: [u8(0x9B), 0x6E] // U+5B3E <cjk>
	`孃`: [u8(0x9B), 0x6F] // U+5B43 <cjk>
	`孅`: [u8(0x9B), 0x70] // U+5B45 <cjk>
	`孀`: [u8(0x9B), 0x71] // U+5B40 <cjk>
	`孑`: [u8(0x9B), 0x72] // U+5B51 <cjk>
	`孕`: [u8(0x9B), 0x73] // U+5B55 <cjk>
	`孚`: [u8(0x9B), 0x74] // U+5B5A <cjk>
	`孛`: [u8(0x9B), 0x75] // U+5B5B <cjk>
	`孥`: [u8(0x9B), 0x76] // U+5B65 <cjk>
	`孩`: [u8(0x9B), 0x77] // U+5B69 <cjk>
	`孰`: [u8(0x9B), 0x78] // U+5B70 <cjk>
	`孳`: [u8(0x9B), 0x79] // U+5B73 <cjk>
	`孵`: [u8(0x9B), 0x7A] // U+5B75 <cjk>
	`學`: [u8(0x9B), 0x7B] // U+5B78 <cjk>
	`斈`: [u8(0x9B), 0x7C] // U+6588 <cjk>
	`孺`: [u8(0x9B), 0x7D] // U+5B7A <cjk>
	`宀`: [u8(0x9B), 0x7E] // U+5B80 <cjk>
	`它`: [u8(0x9B), 0x80] // U+5B83 <cjk>
	`宦`: [u8(0x9B), 0x81] // U+5BA6 <cjk>
	`宸`: [u8(0x9B), 0x82] // U+5BB8 <cjk>
	`寃`: [u8(0x9B), 0x83] // U+5BC3 <cjk>
	`寇`: [u8(0x9B), 0x84] // U+5BC7 <cjk>
	`寉`: [u8(0x9B), 0x85] // U+5BC9 <cjk>
	`寔`: [u8(0x9B), 0x86] // U+5BD4 <cjk>
	`寐`: [u8(0x9B), 0x87] // U+5BD0 <cjk>
	`寤`: [u8(0x9B), 0x88] // U+5BE4 <cjk>
	`實`: [u8(0x9B), 0x89] // U+5BE6 <cjk>
	`寢`: [u8(0x9B), 0x8A] // U+5BE2 <cjk>
	`寞`: [u8(0x9B), 0x8B] // U+5BDE <cjk>
	`寥`: [u8(0x9B), 0x8C] // U+5BE5 <cjk>
	`寫`: [u8(0x9B), 0x8D] // U+5BEB <cjk>
	`寰`: [u8(0x9B), 0x8E] // U+5BF0 <cjk>
	`寶`: [u8(0x9B), 0x8F] // U+5BF6 <cjk>
	`寳`: [u8(0x9B), 0x90] // U+5BF3 <cjk>
	`尅`: [u8(0x9B), 0x91] // U+5C05 <cjk>
	`將`: [u8(0x9B), 0x92] // U+5C07 <cjk>
	`專`: [u8(0x9B), 0x93] // U+5C08 <cjk>
	`對`: [u8(0x9B), 0x94] // U+5C0D <cjk>
	`尓`: [u8(0x9B), 0x95] // U+5C13 <cjk>
	`尠`: [u8(0x9B), 0x96] // U+5C20 <cjk>
	`尢`: [u8(0x9B), 0x97] // U+5C22 <cjk>
	`尨`: [u8(0x9B), 0x98] // U+5C28 <cjk>
	`尸`: [u8(0x9B), 0x99] // U+5C38 <cjk>
	`尹`: [u8(0x9B), 0x9A] // U+5C39 <cjk>
	`屁`: [u8(0x9B), 0x9B] // U+5C41 <cjk>
	`屆`: [u8(0x9B), 0x9C] // U+5C46 <cjk>
	`屎`: [u8(0x9B), 0x9D] // U+5C4E <cjk>
	`屓`: [u8(0x9B), 0x9E] // U+5C53 <cjk>
	`屐`: [u8(0x9B), 0x9F] // U+5C50 <cjk>
	`屏`: [u8(0x9B), 0xA0] // U+5C4F <cjk>
	`孱`: [u8(0x9B), 0xA1] // U+5B71 <cjk>
	`屬`: [u8(0x9B), 0xA2] // U+5C6C <cjk>
	`屮`: [u8(0x9B), 0xA3] // U+5C6E <cjk>
	`乢`: [u8(0x9B), 0xA4] // U+4E62 <cjk>
	`屶`: [u8(0x9B), 0xA5] // U+5C76 <cjk>
	`屹`: [u8(0x9B), 0xA6] // U+5C79 <cjk>
	`岌`: [u8(0x9B), 0xA7] // U+5C8C <cjk>
	`岑`: [u8(0x9B), 0xA8] // U+5C91 <cjk>
	`岔`: [u8(0x9B), 0xA9] // U+5C94 <cjk>
	`妛`: [u8(0x9B), 0xAA] // U+599B <cjk>
	`岫`: [u8(0x9B), 0xAB] // U+5CAB <cjk>
	`岻`: [u8(0x9B), 0xAC] // U+5CBB <cjk>
	`岶`: [u8(0x9B), 0xAD] // U+5CB6 <cjk>
	`岼`: [u8(0x9B), 0xAE] // U+5CBC <cjk>
	`岷`: [u8(0x9B), 0xAF] // U+5CB7 <cjk>
	`峅`: [u8(0x9B), 0xB0] // U+5CC5 <cjk>
	`岾`: [u8(0x9B), 0xB1] // U+5CBE <cjk>
	`峇`: [u8(0x9B), 0xB2] // U+5CC7 <cjk>
	`峙`: [u8(0x9B), 0xB3] // U+5CD9 <cjk>
	`峩`: [u8(0x9B), 0xB4] // U+5CE9 <cjk>
	`峽`: [u8(0x9B), 0xB5] // U+5CFD <cjk>
	`峺`: [u8(0x9B), 0xB6] // U+5CFA <cjk>
	`峭`: [u8(0x9B), 0xB7] // U+5CED <cjk>
	`嶌`: [u8(0x9B), 0xB8] // U+5D8C <cjk>
	`峪`: [u8(0x9B), 0xB9] // U+5CEA <cjk>
	`崋`: [u8(0x9B), 0xBA] // U+5D0B <cjk>
	`崕`: [u8(0x9B), 0xBB] // U+5D15 <cjk>
	`崗`: [u8(0x9B), 0xBC] // U+5D17 <cjk>
	`嵜`: [u8(0x9B), 0xBD] // U+5D5C <cjk>
	`崟`: [u8(0x9B), 0xBE] // U+5D1F <cjk>
	`崛`: [u8(0x9B), 0xBF] // U+5D1B <cjk>
	`崑`: [u8(0x9B), 0xC0] // U+5D11 <cjk>
	`崔`: [u8(0x9B), 0xC1] // U+5D14 <cjk>
	`崢`: [u8(0x9B), 0xC2] // U+5D22 <cjk>
	`崚`: [u8(0x9B), 0xC3] // U+5D1A <cjk>
	`崙`: [u8(0x9B), 0xC4] // U+5D19 <cjk>
	`崘`: [u8(0x9B), 0xC5] // U+5D18 <cjk>
	`嵌`: [u8(0x9B), 0xC6] // U+5D4C <cjk>
	`嵒`: [u8(0x9B), 0xC7] // U+5D52 <cjk>
	`嵎`: [u8(0x9B), 0xC8] // U+5D4E <cjk>
	`嵋`: [u8(0x9B), 0xC9] // U+5D4B <cjk>
	`嵬`: [u8(0x9B), 0xCA] // U+5D6C <cjk>
	`嵳`: [u8(0x9B), 0xCB] // U+5D73 <cjk>
	`嵶`: [u8(0x9B), 0xCC] // U+5D76 <cjk>
	`嶇`: [u8(0x9B), 0xCD] // U+5D87 <cjk>
	`嶄`: [u8(0x9B), 0xCE] // U+5D84 <cjk>
	`嶂`: [u8(0x9B), 0xCF] // U+5D82 <cjk>
	`嶢`: [u8(0x9B), 0xD0] // U+5DA2 <cjk>
	`嶝`: [u8(0x9B), 0xD1] // U+5D9D <cjk>
	`嶬`: [u8(0x9B), 0xD2] // U+5DAC <cjk>
	`嶮`: [u8(0x9B), 0xD3] // U+5DAE <cjk>
	`嶽`: [u8(0x9B), 0xD4] // U+5DBD <cjk>
	`嶐`: [u8(0x9B), 0xD5] // U+5D90 <cjk>
	`嶷`: [u8(0x9B), 0xD6] // U+5DB7 <cjk>
	`嶼`: [u8(0x9B), 0xD7] // U+5DBC <cjk>
	`巉`: [u8(0x9B), 0xD8] // U+5DC9 <cjk>
	`巍`: [u8(0x9B), 0xD9] // U+5DCD <cjk>
	`巓`: [u8(0x9B), 0xDA] // U+5DD3 <cjk>
	`巒`: [u8(0x9B), 0xDB] // U+5DD2 <cjk>
	`巖`: [u8(0x9B), 0xDC] // U+5DD6 <cjk>
	`巛`: [u8(0x9B), 0xDD] // U+5DDB <cjk>
	`巫`: [u8(0x9B), 0xDE] // U+5DEB <cjk>
	`已`: [u8(0x9B), 0xDF] // U+5DF2 <cjk>
	`巵`: [u8(0x9B), 0xE0] // U+5DF5 <cjk>
	`帋`: [u8(0x9B), 0xE1] // U+5E0B <cjk>
	`帚`: [u8(0x9B), 0xE2] // U+5E1A <cjk>
	`帙`: [u8(0x9B), 0xE3] // U+5E19 <cjk>
	`帑`: [u8(0x9B), 0xE4] // U+5E11 <cjk>
	`帛`: [u8(0x9B), 0xE5] // U+5E1B <cjk>
	`帶`: [u8(0x9B), 0xE6] // U+5E36 <cjk>
	`帷`: [u8(0x9B), 0xE7] // U+5E37 <cjk>
	`幄`: [u8(0x9B), 0xE8] // U+5E44 <cjk>
	`幃`: [u8(0x9B), 0xE9] // U+5E43 <cjk>
	`幀`: [u8(0x9B), 0xEA] // U+5E40 <cjk>
	`幎`: [u8(0x9B), 0xEB] // U+5E4E <cjk>
	`幗`: [u8(0x9B), 0xEC] // U+5E57 <cjk>
	`幔`: [u8(0x9B), 0xED] // U+5E54 <cjk>
	`幟`: [u8(0x9B), 0xEE] // U+5E5F <cjk>
	`幢`: [u8(0x9B), 0xEF] // U+5E62 <cjk>
	`幤`: [u8(0x9B), 0xF0] // U+5E64 <cjk>
	`幇`: [u8(0x9B), 0xF1] // U+5E47 <cjk>
	`幵`: [u8(0x9B), 0xF2] // U+5E75 <cjk>
	`并`: [u8(0x9B), 0xF3] // U+5E76 <cjk>
	`幺`: [u8(0x9B), 0xF4] // U+5E7A <cjk>
	`麼`: [u8(0x9B), 0xF5] // U+9EBC <cjk>
	`广`: [u8(0x9B), 0xF6] // U+5E7F <cjk>
	`庠`: [u8(0x9B), 0xF7] // U+5EA0 <cjk>
	`廁`: [u8(0x9B), 0xF8] // U+5EC1 <cjk>
	`廂`: [u8(0x9B), 0xF9] // U+5EC2 <cjk>
	`廈`: [u8(0x9B), 0xFA] // U+5EC8 <cjk>
	`廐`: [u8(0x9B), 0xFB] // U+5ED0 <cjk>
	`廏`: [u8(0x9B), 0xFC] // U+5ECF <cjk>
	`廖`: [u8(0x9C), 0x40] // U+5ED6 <cjk>
	`廣`: [u8(0x9C), 0x41] // U+5EE3 <cjk>
	`廝`: [u8(0x9C), 0x42] // U+5EDD <cjk>
	`廚`: [u8(0x9C), 0x43] // U+5EDA <cjk>
	`廛`: [u8(0x9C), 0x44] // U+5EDB <cjk>
	`廢`: [u8(0x9C), 0x45] // U+5EE2 <cjk>
	`廡`: [u8(0x9C), 0x46] // U+5EE1 <cjk>
	`廨`: [u8(0x9C), 0x47] // U+5EE8 <cjk>
	`廩`: [u8(0x9C), 0x48] // U+5EE9 <cjk>
	`廬`: [u8(0x9C), 0x49] // U+5EEC <cjk>
	`廱`: [u8(0x9C), 0x4A] // U+5EF1 <cjk>
	`廳`: [u8(0x9C), 0x4B] // U+5EF3 <cjk>
	`廰`: [u8(0x9C), 0x4C] // U+5EF0 <cjk>
	`廴`: [u8(0x9C), 0x4D] // U+5EF4 <cjk>
	`廸`: [u8(0x9C), 0x4E] // U+5EF8 <cjk>
	`廾`: [u8(0x9C), 0x4F] // U+5EFE <cjk>
	`弃`: [u8(0x9C), 0x50] // U+5F03 <cjk>
	`弉`: [u8(0x9C), 0x51] // U+5F09 <cjk>
	`彝`: [u8(0x9C), 0x52] // U+5F5D <cjk>
	`彜`: [u8(0x9C), 0x53] // U+5F5C <cjk>
	`弋`: [u8(0x9C), 0x54] // U+5F0B <cjk>
	`弑`: [u8(0x9C), 0x55] // U+5F11 <cjk>
	`弖`: [u8(0x9C), 0x56] // U+5F16 <cjk>
	`弩`: [u8(0x9C), 0x57] // U+5F29 <cjk>
	`弭`: [u8(0x9C), 0x58] // U+5F2D <cjk>
	`弸`: [u8(0x9C), 0x59] // U+5F38 <cjk>
	`彁`: [u8(0x9C), 0x5A] // U+5F41 <cjk>
	`彈`: [u8(0x9C), 0x5B] // U+5F48 <cjk>
	`彌`: [u8(0x9C), 0x5C] // U+5F4C <cjk>
	`彎`: [u8(0x9C), 0x5D] // U+5F4E <cjk>
	`弯`: [u8(0x9C), 0x5E] // U+5F2F <cjk>
	`彑`: [u8(0x9C), 0x5F] // U+5F51 <cjk>
	`彖`: [u8(0x9C), 0x60] // U+5F56 <cjk>
	`彗`: [u8(0x9C), 0x61] // U+5F57 <cjk>
	`彙`: [u8(0x9C), 0x62] // U+5F59 <cjk>
	`彡`: [u8(0x9C), 0x63] // U+5F61 <cjk>
	`彭`: [u8(0x9C), 0x64] // U+5F6D <cjk>
	`彳`: [u8(0x9C), 0x65] // U+5F73 <cjk>
	`彷`: [u8(0x9C), 0x66] // U+5F77 <cjk>
	`徃`: [u8(0x9C), 0x67] // U+5F83 <cjk>
	`徂`: [u8(0x9C), 0x68] // U+5F82 <cjk>
	`彿`: [u8(0x9C), 0x69] // U+5F7F <cjk>
	`徊`: [u8(0x9C), 0x6A] // U+5F8A <cjk>
	`很`: [u8(0x9C), 0x6B] // U+5F88 <cjk>
	`徑`: [u8(0x9C), 0x6C] // U+5F91 <cjk>
	`徇`: [u8(0x9C), 0x6D] // U+5F87 <cjk>
	`從`: [u8(0x9C), 0x6E] // U+5F9E <cjk>
	`徙`: [u8(0x9C), 0x6F] // U+5F99 <cjk>
	`徘`: [u8(0x9C), 0x70] // U+5F98 <cjk>
	`徠`: [u8(0x9C), 0x71] // U+5FA0 <cjk>
	`徨`: [u8(0x9C), 0x72] // U+5FA8 <cjk>
	`徭`: [u8(0x9C), 0x73] // U+5FAD <cjk>
	`徼`: [u8(0x9C), 0x74] // U+5FBC <cjk>
	`忖`: [u8(0x9C), 0x75] // U+5FD6 <cjk>
	`忻`: [u8(0x9C), 0x76] // U+5FFB <cjk>
	`忤`: [u8(0x9C), 0x77] // U+5FE4 <cjk>
	`忸`: [u8(0x9C), 0x78] // U+5FF8 <cjk>
	`忱`: [u8(0x9C), 0x79] // U+5FF1 <cjk>
	`忝`: [u8(0x9C), 0x7A] // U+5FDD <cjk>
	`悳`: [u8(0x9C), 0x7B] // U+60B3 <cjk>
	`忿`: [u8(0x9C), 0x7C] // U+5FFF <cjk>
	`怡`: [u8(0x9C), 0x7D] // U+6021 <cjk>
	`恠`: [u8(0x9C), 0x7E] // U+6060 <cjk>
	`怙`: [u8(0x9C), 0x80] // U+6019 <cjk>
	`怐`: [u8(0x9C), 0x81] // U+6010 <cjk>
	`怩`: [u8(0x9C), 0x82] // U+6029 <cjk>
	`怎`: [u8(0x9C), 0x83] // U+600E <cjk>
	`怱`: [u8(0x9C), 0x84] // U+6031 <cjk>
	`怛`: [u8(0x9C), 0x85] // U+601B <cjk>
	`怕`: [u8(0x9C), 0x86] // U+6015 <cjk>
	`怫`: [u8(0x9C), 0x87] // U+602B <cjk>
	`怦`: [u8(0x9C), 0x88] // U+6026 <cjk>
	`怏`: [u8(0x9C), 0x89] // U+600F <cjk>
	`怺`: [u8(0x9C), 0x8A] // U+603A <cjk>
	`恚`: [u8(0x9C), 0x8B] // U+605A <cjk>
	`恁`: [u8(0x9C), 0x8C] // U+6041 <cjk>
	`恪`: [u8(0x9C), 0x8D] // U+606A <cjk>
	`恷`: [u8(0x9C), 0x8E] // U+6077 <cjk>
	`恟`: [u8(0x9C), 0x8F] // U+605F <cjk>
	`恊`: [u8(0x9C), 0x90] // U+604A <cjk>
	`恆`: [u8(0x9C), 0x91] // U+6046 <cjk>
	`恍`: [u8(0x9C), 0x92] // U+604D <cjk>
	`恣`: [u8(0x9C), 0x93] // U+6063 <cjk>
	`恃`: [u8(0x9C), 0x94] // U+6043 <cjk>
	`恤`: [u8(0x9C), 0x95] // U+6064 <cjk>
	`恂`: [u8(0x9C), 0x96] // U+6042 <cjk>
	`恬`: [u8(0x9C), 0x97] // U+606C <cjk>
	`恫`: [u8(0x9C), 0x98] // U+606B <cjk>
	`恙`: [u8(0x9C), 0x99] // U+6059 <cjk>
	`悁`: [u8(0x9C), 0x9A] // U+6081 <cjk>
	`悍`: [u8(0x9C), 0x9B] // U+608D <cjk>
	`惧`: [u8(0x9C), 0x9C] // U+60E7 <cjk>
	`悃`: [u8(0x9C), 0x9D] // U+6083 <cjk>
	`悚`: [u8(0x9C), 0x9E] // U+609A <cjk>
	`悄`: [u8(0x9C), 0x9F] // U+6084 <cjk>
	`悛`: [u8(0x9C), 0xA0] // U+609B <cjk>
	`悖`: [u8(0x9C), 0xA1] // U+6096 <cjk>
	`悗`: [u8(0x9C), 0xA2] // U+6097 <cjk>
	`悒`: [u8(0x9C), 0xA3] // U+6092 <cjk>
	`悧`: [u8(0x9C), 0xA4] // U+60A7 <cjk>
	`悋`: [u8(0x9C), 0xA5] // U+608B <cjk>
	`惡`: [u8(0x9C), 0xA6] // U+60E1 <cjk>
	`悸`: [u8(0x9C), 0xA7] // U+60B8 <cjk>
	`惠`: [u8(0x9C), 0xA8] // U+60E0 <cjk>
	`惓`: [u8(0x9C), 0xA9] // U+60D3 <cjk>
	`悴`: [u8(0x9C), 0xAA] // U+60B4 <cjk>
	`忰`: [u8(0x9C), 0xAB] // U+5FF0 <cjk>
	`悽`: [u8(0x9C), 0xAC] // U+60BD <cjk>
	`惆`: [u8(0x9C), 0xAD] // U+60C6 <cjk>
	`悵`: [u8(0x9C), 0xAE] // U+60B5 <cjk>
	`惘`: [u8(0x9C), 0xAF] // U+60D8 <cjk>
	`慍`: [u8(0x9C), 0xB0] // U+614D <cjk>
	`愕`: [u8(0x9C), 0xB1] // U+6115 <cjk>
	`愆`: [u8(0x9C), 0xB2] // U+6106 <cjk>
	`惶`: [u8(0x9C), 0xB3] // U+60F6 <cjk>
	`惷`: [u8(0x9C), 0xB4] // U+60F7 <cjk>
	`愀`: [u8(0x9C), 0xB5] // U+6100 <cjk>
	`惴`: [u8(0x9C), 0xB6] // U+60F4 <cjk>
	`惺`: [u8(0x9C), 0xB7] // U+60FA <cjk>
	`愃`: [u8(0x9C), 0xB8] // U+6103 <cjk>
	`愡`: [u8(0x9C), 0xB9] // U+6121 <cjk>
	`惻`: [u8(0x9C), 0xBA] // U+60FB <cjk>
	`惱`: [u8(0x9C), 0xBB] // U+60F1 <cjk>
	`愍`: [u8(0x9C), 0xBC] // U+610D <cjk>
	`愎`: [u8(0x9C), 0xBD] // U+610E <cjk>
	`慇`: [u8(0x9C), 0xBE] // U+6147 <cjk>
	`愾`: [u8(0x9C), 0xBF] // U+613E <cjk>
	`愨`: [u8(0x9C), 0xC0] // U+6128 <cjk>
	`愧`: [u8(0x9C), 0xC1] // U+6127 <cjk>
	`慊`: [u8(0x9C), 0xC2] // U+614A <cjk>
	`愿`: [u8(0x9C), 0xC3] // U+613F <cjk>
	`愼`: [u8(0x9C), 0xC4] // U+613C <cjk>
	`愬`: [u8(0x9C), 0xC5] // U+612C <cjk>
	`愴`: [u8(0x9C), 0xC6] // U+6134 <cjk>
	`愽`: [u8(0x9C), 0xC7] // U+613D <cjk>
	`慂`: [u8(0x9C), 0xC8] // U+6142 <cjk>
	`慄`: [u8(0x9C), 0xC9] // U+6144 <cjk>
	`慳`: [u8(0x9C), 0xCA] // U+6173 <cjk>
	`慷`: [u8(0x9C), 0xCB] // U+6177 <cjk>
	`慘`: [u8(0x9C), 0xCC] // U+6158 <cjk>
	`慙`: [u8(0x9C), 0xCD] // U+6159 <cjk>
	`慚`: [u8(0x9C), 0xCE] // U+615A <cjk>
	`慫`: [u8(0x9C), 0xCF] // U+616B <cjk>
	`慴`: [u8(0x9C), 0xD0] // U+6174 <cjk>
	`慯`: [u8(0x9C), 0xD1] // U+616F <cjk>
	`慥`: [u8(0x9C), 0xD2] // U+6165 <cjk>
	`慱`: [u8(0x9C), 0xD3] // U+6171 <cjk>
	`慟`: [u8(0x9C), 0xD4] // U+615F <cjk>
	`慝`: [u8(0x9C), 0xD5] // U+615D <cjk>
	`慓`: [u8(0x9C), 0xD6] // U+6153 <cjk>
	`慵`: [u8(0x9C), 0xD7] // U+6175 <cjk>
	`憙`: [u8(0x9C), 0xD8] // U+6199 <cjk>
	`憖`: [u8(0x9C), 0xD9] // U+6196 <cjk>
	`憇`: [u8(0x9C), 0xDA] // U+6187 <cjk>
	`憬`: [u8(0x9C), 0xDB] // U+61AC <cjk>
	`憔`: [u8(0x9C), 0xDC] // U+6194 <cjk>
	`憚`: [u8(0x9C), 0xDD] // U+619A <cjk>
	`憊`: [u8(0x9C), 0xDE] // U+618A <cjk>
	`憑`: [u8(0x9C), 0xDF] // U+6191 <cjk>
	`憫`: [u8(0x9C), 0xE0] // U+61AB <cjk>
	`憮`: [u8(0x9C), 0xE1] // U+61AE <cjk>
	`懌`: [u8(0x9C), 0xE2] // U+61CC <cjk>
	`懊`: [u8(0x9C), 0xE3] // U+61CA <cjk>
	`應`: [u8(0x9C), 0xE4] // U+61C9 <cjk>
	`懷`: [u8(0x9C), 0xE5] // U+61F7 <cjk>
	`懈`: [u8(0x9C), 0xE6] // U+61C8 <cjk>
	`懃`: [u8(0x9C), 0xE7] // U+61C3 <cjk>
	`懆`: [u8(0x9C), 0xE8] // U+61C6 <cjk>
	`憺`: [u8(0x9C), 0xE9] // U+61BA <cjk>
	`懋`: [u8(0x9C), 0xEA] // U+61CB <cjk>
	`罹`: [u8(0x9C), 0xEB] // U+7F79 <cjk>
	`懍`: [u8(0x9C), 0xEC] // U+61CD <cjk>
	`懦`: [u8(0x9C), 0xED] // U+61E6 <cjk>
	`懣`: [u8(0x9C), 0xEE] // U+61E3 <cjk>
	`懶`: [u8(0x9C), 0xEF] // U+61F6 <cjk>
	`懺`: [u8(0x9C), 0xF0] // U+61FA <cjk>
	`懴`: [u8(0x9C), 0xF1] // U+61F4 <cjk>
	`懿`: [u8(0x9C), 0xF2] // U+61FF <cjk>
	`懽`: [u8(0x9C), 0xF3] // U+61FD <cjk>
	`懼`: [u8(0x9C), 0xF4] // U+61FC <cjk>
	`懾`: [u8(0x9C), 0xF5] // U+61FE <cjk>
	`戀`: [u8(0x9C), 0xF6] // U+6200 <cjk>
	`戈`: [u8(0x9C), 0xF7] // U+6208 <cjk>
	`戉`: [u8(0x9C), 0xF8] // U+6209 <cjk>
	`戍`: [u8(0x9C), 0xF9] // U+620D <cjk>
	`戌`: [u8(0x9C), 0xFA] // U+620C <cjk>
	`戔`: [u8(0x9C), 0xFB] // U+6214 <cjk>
	`戛`: [u8(0x9C), 0xFC] // U+621B <cjk>
	`戞`: [u8(0x9D), 0x40] // U+621E <cjk>
	`戡`: [u8(0x9D), 0x41] // U+6221 <cjk>
	`截`: [u8(0x9D), 0x42] // U+622A <cjk>
	`戮`: [u8(0x9D), 0x43] // U+622E <cjk>
	`戰`: [u8(0x9D), 0x44] // U+6230 <cjk>
	`戲`: [u8(0x9D), 0x45] // U+6232 <cjk>
	`戳`: [u8(0x9D), 0x46] // U+6233 <cjk>
	`扁`: [u8(0x9D), 0x47] // U+6241 <cjk>
	`扎`: [u8(0x9D), 0x48] // U+624E <cjk>
	`扞`: [u8(0x9D), 0x49] // U+625E <cjk>
	`扣`: [u8(0x9D), 0x4A] // U+6263 <cjk>
	`扛`: [u8(0x9D), 0x4B] // U+625B <cjk>
	`扠`: [u8(0x9D), 0x4C] // U+6260 <cjk>
	`扨`: [u8(0x9D), 0x4D] // U+6268 <cjk>
	`扼`: [u8(0x9D), 0x4E] // U+627C <cjk>
	`抂`: [u8(0x9D), 0x4F] // U+6282 <cjk>
	`抉`: [u8(0x9D), 0x50] // U+6289 <cjk>
	`找`: [u8(0x9D), 0x51] // U+627E <cjk>
	`抒`: [u8(0x9D), 0x52] // U+6292 <cjk>
	`抓`: [u8(0x9D), 0x53] // U+6293 <cjk>
	`抖`: [u8(0x9D), 0x54] // U+6296 <cjk>
	`拔`: [u8(0x9D), 0x55] // U+62D4 <cjk>
	`抃`: [u8(0x9D), 0x56] // U+6283 <cjk>
	`抔`: [u8(0x9D), 0x57] // U+6294 <cjk>
	`拗`: [u8(0x9D), 0x58] // U+62D7 <cjk>
	`拑`: [u8(0x9D), 0x59] // U+62D1 <cjk>
	`抻`: [u8(0x9D), 0x5A] // U+62BB <cjk>
	`拏`: [u8(0x9D), 0x5B] // U+62CF <cjk>
	`拿`: [u8(0x9D), 0x5C] // U+62FF <cjk>
	`拆`: [u8(0x9D), 0x5D] // U+62C6 <cjk>
	`擔`: [u8(0x9D), 0x5E] // U+64D4 <cjk>
	`拈`: [u8(0x9D), 0x5F] // U+62C8 <cjk>
	`拜`: [u8(0x9D), 0x60] // U+62DC <cjk>
	`拌`: [u8(0x9D), 0x61] // U+62CC <cjk>
	`拊`: [u8(0x9D), 0x62] // U+62CA <cjk>
	`拂`: [u8(0x9D), 0x63] // U+62C2 <cjk>
	`拇`: [u8(0x9D), 0x64] // U+62C7 <cjk>
	`抛`: [u8(0x9D), 0x65] // U+629B <cjk>
	`拉`: [u8(0x9D), 0x66] // U+62C9 <cjk>
	`挌`: [u8(0x9D), 0x67] // U+630C <cjk>
	`拮`: [u8(0x9D), 0x68] // U+62EE <cjk>
	`拱`: [u8(0x9D), 0x69] // U+62F1 <cjk>
	`挧`: [u8(0x9D), 0x6A] // U+6327 <cjk>
	`挂`: [u8(0x9D), 0x6B] // U+6302 <cjk>
	`挈`: [u8(0x9D), 0x6C] // U+6308 <cjk>
	`拯`: [u8(0x9D), 0x6D] // U+62EF <cjk>
	`拵`: [u8(0x9D), 0x6E] // U+62F5 <cjk>
	`捐`: [u8(0x9D), 0x6F] // U+6350 <cjk>
	`挾`: [u8(0x9D), 0x70] // U+633E <cjk>
	`捍`: [u8(0x9D), 0x71] // U+634D <cjk>
	`搜`: [u8(0x9D), 0x72] // U+641C <cjk>
	`捏`: [u8(0x9D), 0x73] // U+634F <cjk>
	`掖`: [u8(0x9D), 0x74] // U+6396 <cjk>
	`掎`: [u8(0x9D), 0x75] // U+638E <cjk>
	`掀`: [u8(0x9D), 0x76] // U+6380 <cjk>
	`掫`: [u8(0x9D), 0x77] // U+63AB <cjk>
	`捶`: [u8(0x9D), 0x78] // U+6376 <cjk>
	`掣`: [u8(0x9D), 0x79] // U+63A3 <cjk>
	`掏`: [u8(0x9D), 0x7A] // U+638F <cjk>
	`掉`: [u8(0x9D), 0x7B] // U+6389 <cjk>
	`掟`: [u8(0x9D), 0x7C] // U+639F <cjk>
	`掵`: [u8(0x9D), 0x7D] // U+63B5 <cjk>
	`捫`: [u8(0x9D), 0x7E] // U+636B <cjk>
	`捩`: [u8(0x9D), 0x80] // U+6369 <cjk>
	`掾`: [u8(0x9D), 0x81] // U+63BE <cjk>
	`揩`: [u8(0x9D), 0x82] // U+63E9 <cjk>
	`揀`: [u8(0x9D), 0x83] // U+63C0 <cjk>
	`揆`: [u8(0x9D), 0x84] // U+63C6 <cjk>
	`揣`: [u8(0x9D), 0x85] // U+63E3 <cjk>
	`揉`: [u8(0x9D), 0x86] // U+63C9 <cjk>
	`插`: [u8(0x9D), 0x87] // U+63D2 <cjk>
	`揶`: [u8(0x9D), 0x88] // U+63F6 <cjk>
	`揄`: [u8(0x9D), 0x89] // U+63C4 <cjk>
	`搖`: [u8(0x9D), 0x8A] // U+6416 <cjk>
	`搴`: [u8(0x9D), 0x8B] // U+6434 <cjk>
	`搆`: [u8(0x9D), 0x8C] // U+6406 <cjk>
	`搓`: [u8(0x9D), 0x8D] // U+6413 <cjk>
	`搦`: [u8(0x9D), 0x8E] // U+6426 <cjk>
	`搶`: [u8(0x9D), 0x8F] // U+6436 <cjk>
	`攝`: [u8(0x9D), 0x90] // U+651D <cjk>
	`搗`: [u8(0x9D), 0x91] // U+6417 <cjk>
	`搨`: [u8(0x9D), 0x92] // U+6428 <cjk>
	`搏`: [u8(0x9D), 0x93] // U+640F <cjk>
	`摧`: [u8(0x9D), 0x94] // U+6467 <cjk>
	`摯`: [u8(0x9D), 0x95] // U+646F <cjk>
	`摶`: [u8(0x9D), 0x96] // U+6476 <cjk>
	`摎`: [u8(0x9D), 0x97] // U+644E <cjk>
	`攪`: [u8(0x9D), 0x98] // U+652A <cjk>
	`撕`: [u8(0x9D), 0x99] // U+6495 <cjk>
	`撓`: [u8(0x9D), 0x9A] // U+6493 <cjk>
	`撥`: [u8(0x9D), 0x9B] // U+64A5 <cjk>
	`撩`: [u8(0x9D), 0x9C] // U+64A9 <cjk>
	`撈`: [u8(0x9D), 0x9D] // U+6488 <cjk>
	`撼`: [u8(0x9D), 0x9E] // U+64BC <cjk>
	`據`: [u8(0x9D), 0x9F] // U+64DA <cjk>
	`擒`: [u8(0x9D), 0xA0] // U+64D2 <cjk>
	`擅`: [u8(0x9D), 0xA1] // U+64C5 <cjk>
	`擇`: [u8(0x9D), 0xA2] // U+64C7 <cjk>
	`撻`: [u8(0x9D), 0xA3] // U+64BB <cjk>
	`擘`: [u8(0x9D), 0xA4] // U+64D8 <cjk>
	`擂`: [u8(0x9D), 0xA5] // U+64C2 <cjk>
	`擱`: [u8(0x9D), 0xA6] // U+64F1 <cjk>
	`擧`: [u8(0x9D), 0xA7] // U+64E7 <cjk>
	`舉`: [u8(0x9D), 0xA8] // U+8209 <cjk>
	`擠`: [u8(0x9D), 0xA9] // U+64E0 <cjk>
	`擡`: [u8(0x9D), 0xAA] // U+64E1 <cjk>
	`抬`: [u8(0x9D), 0xAB] // U+62AC <cjk>
	`擣`: [u8(0x9D), 0xAC] // U+64E3 <cjk>
	`擯`: [u8(0x9D), 0xAD] // U+64EF <cjk>
	`攬`: [u8(0x9D), 0xAE] // U+652C <cjk>
	`擶`: [u8(0x9D), 0xAF] // U+64F6 <cjk>
	`擴`: [u8(0x9D), 0xB0] // U+64F4 <cjk>
	`擲`: [u8(0x9D), 0xB1] // U+64F2 <cjk>
	`擺`: [u8(0x9D), 0xB2] // U+64FA <cjk>
	`攀`: [u8(0x9D), 0xB3] // U+6500 <cjk>
	`擽`: [u8(0x9D), 0xB4] // U+64FD <cjk>
	`攘`: [u8(0x9D), 0xB5] // U+6518 <cjk>
	`攜`: [u8(0x9D), 0xB6] // U+651C <cjk>
	`攅`: [u8(0x9D), 0xB7] // U+6505 <cjk>
	`攤`: [u8(0x9D), 0xB8] // U+6524 <cjk>
	`攣`: [u8(0x9D), 0xB9] // U+6523 <cjk>
	`攫`: [u8(0x9D), 0xBA] // U+652B <cjk>
	`攴`: [u8(0x9D), 0xBB] // U+6534 <cjk>
	`攵`: [u8(0x9D), 0xBC] // U+6535 <cjk>
	`攷`: [u8(0x9D), 0xBD] // U+6537 <cjk>
	`收`: [u8(0x9D), 0xBE] // U+6536 <cjk>
	`攸`: [u8(0x9D), 0xBF] // U+6538 <cjk>
	`畋`: [u8(0x9D), 0xC0] // U+754B <cjk>
	`效`: [u8(0x9D), 0xC1] // U+6548 <cjk>
	`敖`: [u8(0x9D), 0xC2] // U+6556 <cjk>
	`敕`: [u8(0x9D), 0xC3] // U+6555 <cjk>
	`敍`: [u8(0x9D), 0xC4] // U+654D <cjk>
	`敘`: [u8(0x9D), 0xC5] // U+6558 <cjk>
	`敞`: [u8(0x9D), 0xC6] // U+655E <cjk>
	`敝`: [u8(0x9D), 0xC7] // U+655D <cjk>
	`敲`: [u8(0x9D), 0xC8] // U+6572 <cjk>
	`數`: [u8(0x9D), 0xC9] // U+6578 <cjk>
	`斂`: [u8(0x9D), 0xCA] // U+6582 <cjk>
	`斃`: [u8(0x9D), 0xCB] // U+6583 <cjk>
	`變`: [u8(0x9D), 0xCC] // U+8B8A <cjk>
	`斛`: [u8(0x9D), 0xCD] // U+659B <cjk>
	`斟`: [u8(0x9D), 0xCE] // U+659F <cjk>
	`斫`: [u8(0x9D), 0xCF] // U+65AB <cjk>
	`斷`: [u8(0x9D), 0xD0] // U+65B7 <cjk>
	`旃`: [u8(0x9D), 0xD1] // U+65C3 <cjk>
	`旆`: [u8(0x9D), 0xD2] // U+65C6 <cjk>
	`旁`: [u8(0x9D), 0xD3] // U+65C1 <cjk>
	`旄`: [u8(0x9D), 0xD4] // U+65C4 <cjk>
	`旌`: [u8(0x9D), 0xD5] // U+65CC <cjk>
	`旒`: [u8(0x9D), 0xD6] // U+65D2 <cjk>
	`旛`: [u8(0x9D), 0xD7] // U+65DB <cjk>
	`旙`: [u8(0x9D), 0xD8] // U+65D9 <cjk>
	`无`: [u8(0x9D), 0xD9] // U+65E0 <cjk>
	`旡`: [u8(0x9D), 0xDA] // U+65E1 <cjk>
	`旱`: [u8(0x9D), 0xDB] // U+65F1 <cjk>
	`杲`: [u8(0x9D), 0xDC] // U+6772 <cjk>
	`昊`: [u8(0x9D), 0xDD] // U+660A <cjk>
	`昃`: [u8(0x9D), 0xDE] // U+6603 <cjk>
	`旻`: [u8(0x9D), 0xDF] // U+65FB <cjk>
	`杳`: [u8(0x9D), 0xE0] // U+6773 <cjk>
	`昵`: [u8(0x9D), 0xE1] // U+6635 <cjk>
	`昶`: [u8(0x9D), 0xE2] // U+6636 <cjk>
	`昴`: [u8(0x9D), 0xE3] // U+6634 <cjk>
	`昜`: [u8(0x9D), 0xE4] // U+661C <cjk>
	`晏`: [u8(0x9D), 0xE5] // U+664F <cjk>
	`晄`: [u8(0x9D), 0xE6] // U+6644 <cjk>
	`晉`: [u8(0x9D), 0xE7] // U+6649 <cjk>
	`晁`: [u8(0x9D), 0xE8] // U+6641 <cjk>
	`晞`: [u8(0x9D), 0xE9] // U+665E <cjk>
	`晝`: [u8(0x9D), 0xEA] // U+665D <cjk>
	`晤`: [u8(0x9D), 0xEB] // U+6664 <cjk>
	`晧`: [u8(0x9D), 0xEC] // U+6667 <cjk>
	`晨`: [u8(0x9D), 0xED] // U+6668 <cjk>
	`晟`: [u8(0x9D), 0xEE] // U+665F <cjk>
	`晢`: [u8(0x9D), 0xEF] // U+6662 <cjk>
	`晰`: [u8(0x9D), 0xF0] // U+6670 <cjk>
	`暃`: [u8(0x9D), 0xF1] // U+6683 <cjk>
	`暈`: [u8(0x9D), 0xF2] // U+6688 <cjk>
	`暎`: [u8(0x9D), 0xF3] // U+668E <cjk>
	`暉`: [u8(0x9D), 0xF4] // U+6689 <cjk>
	`暄`: [u8(0x9D), 0xF5] // U+6684 <cjk>
	`暘`: [u8(0x9D), 0xF6] // U+6698 <cjk>
	`暝`: [u8(0x9D), 0xF7] // U+669D <cjk>
	`曁`: [u8(0x9D), 0xF8] // U+66C1 <cjk>
	`暹`: [u8(0x9D), 0xF9] // U+66B9 <cjk>
	`曉`: [u8(0x9D), 0xFA] // U+66C9 <cjk>
	`暾`: [u8(0x9D), 0xFB] // U+66BE <cjk>
	`暼`: [u8(0x9D), 0xFC] // U+66BC <cjk>
	`曄`: [u8(0x9E), 0x40] // U+66C4 <cjk>
	`暸`: [u8(0x9E), 0x41] // U+66B8 <cjk>
	`曖`: [u8(0x9E), 0x42] // U+66D6 <cjk>
	`曚`: [u8(0x9E), 0x43] // U+66DA <cjk>
	`曠`: [u8(0x9E), 0x44] // U+66E0 <cjk>
	`昿`: [u8(0x9E), 0x45] // U+663F <cjk>
	`曦`: [u8(0x9E), 0x46] // U+66E6 <cjk>
	`曩`: [u8(0x9E), 0x47] // U+66E9 <cjk>
	`曰`: [u8(0x9E), 0x48] // U+66F0 <cjk>
	`曵`: [u8(0x9E), 0x49] // U+66F5 <cjk>
	`曷`: [u8(0x9E), 0x4A] // U+66F7 <cjk>
	`朏`: [u8(0x9E), 0x4B] // U+670F <cjk>
	`朖`: [u8(0x9E), 0x4C] // U+6716 <cjk>
	`朞`: [u8(0x9E), 0x4D] // U+671E <cjk>
	`朦`: [u8(0x9E), 0x4E] // U+6726 <cjk>
	`朧`: [u8(0x9E), 0x4F] // U+6727 <cjk>
	`霸`: [u8(0x9E), 0x50] // U+9738 <cjk>
	`朮`: [u8(0x9E), 0x51] // U+672E <cjk>
	`朿`: [u8(0x9E), 0x52] // U+673F <cjk>
	`朶`: [u8(0x9E), 0x53] // U+6736 <cjk>
	`杁`: [u8(0x9E), 0x54] // U+6741 <cjk>
	`朸`: [u8(0x9E), 0x55] // U+6738 <cjk>
	`朷`: [u8(0x9E), 0x56] // U+6737 <cjk>
	`杆`: [u8(0x9E), 0x57] // U+6746 <cjk>
	`杞`: [u8(0x9E), 0x58] // U+675E <cjk>
	`杠`: [u8(0x9E), 0x59] // U+6760 <cjk>
	`杙`: [u8(0x9E), 0x5A] // U+6759 <cjk>
	`杣`: [u8(0x9E), 0x5B] // U+6763 <cjk>
	`杤`: [u8(0x9E), 0x5C] // U+6764 <cjk>
	`枉`: [u8(0x9E), 0x5D] // U+6789 <cjk>
	`杰`: [u8(0x9E), 0x5E] // U+6770 <cjk>
	`枩`: [u8(0x9E), 0x5F] // U+67A9 <cjk>
	`杼`: [u8(0x9E), 0x60] // U+677C <cjk>
	`杪`: [u8(0x9E), 0x61] // U+676A <cjk>
	`枌`: [u8(0x9E), 0x62] // U+678C <cjk>
	`枋`: [u8(0x9E), 0x63] // U+678B <cjk>
	`枦`: [u8(0x9E), 0x64] // U+67A6 <cjk>
	`枡`: [u8(0x9E), 0x65] // U+67A1 <cjk>
	`枅`: [u8(0x9E), 0x66] // U+6785 <cjk>
	`枷`: [u8(0x9E), 0x67] // U+67B7 <cjk>
	`柯`: [u8(0x9E), 0x68] // U+67EF <cjk>
	`枴`: [u8(0x9E), 0x69] // U+67B4 <cjk>
	`柬`: [u8(0x9E), 0x6A] // U+67EC <cjk>
	`枳`: [u8(0x9E), 0x6B] // U+67B3 <cjk>
	`柩`: [u8(0x9E), 0x6C] // U+67E9 <cjk>
	`枸`: [u8(0x9E), 0x6D] // U+67B8 <cjk>
	`柤`: [u8(0x9E), 0x6E] // U+67E4 <cjk>
	`柞`: [u8(0x9E), 0x6F] // U+67DE <cjk>
	`柝`: [u8(0x9E), 0x70] // U+67DD <cjk>
	`柢`: [u8(0x9E), 0x71] // U+67E2 <cjk>
	`柮`: [u8(0x9E), 0x72] // U+67EE <cjk>
	`枹`: [u8(0x9E), 0x73] // U+67B9 <cjk>
	`柎`: [u8(0x9E), 0x74] // U+67CE <cjk>
	`柆`: [u8(0x9E), 0x75] // U+67C6 <cjk>
	`柧`: [u8(0x9E), 0x76] // U+67E7 <cjk>
	`檜`: [u8(0x9E), 0x77] // U+6A9C <cjk>
	`栞`: [u8(0x9E), 0x78] // U+681E <cjk>
	`框`: [u8(0x9E), 0x79] // U+6846 <cjk>
	`栩`: [u8(0x9E), 0x7A] // U+6829 <cjk>
	`桀`: [u8(0x9E), 0x7B] // U+6840 <cjk>
	`桍`: [u8(0x9E), 0x7C] // U+684D <cjk>
	`栲`: [u8(0x9E), 0x7D] // U+6832 <cjk>
	`桎`: [u8(0x9E), 0x7E] // U+684E <cjk>
	`梳`: [u8(0x9E), 0x80] // U+68B3 <cjk>
	`栫`: [u8(0x9E), 0x81] // U+682B <cjk>
	`桙`: [u8(0x9E), 0x82] // U+6859 <cjk>
	`档`: [u8(0x9E), 0x83] // U+6863 <cjk>
	`桷`: [u8(0x9E), 0x84] // U+6877 <cjk>
	`桿`: [u8(0x9E), 0x85] // U+687F <cjk>
	`梟`: [u8(0x9E), 0x86] // U+689F <cjk>
	`梏`: [u8(0x9E), 0x87] // U+688F <cjk>
	`梭`: [u8(0x9E), 0x88] // U+68AD <cjk>
	`梔`: [u8(0x9E), 0x89] // U+6894 <cjk>
	`條`: [u8(0x9E), 0x8A] // U+689D <cjk>
	`梛`: [u8(0x9E), 0x8B] // U+689B <cjk>
	`梃`: [u8(0x9E), 0x8C] // U+6883 <cjk>
	`檮`: [u8(0x9E), 0x8D] // U+6AAE <cjk>
	`梹`: [u8(0x9E), 0x8E] // U+68B9 <cjk>
	`桴`: [u8(0x9E), 0x8F] // U+6874 <cjk>
	`梵`: [u8(0x9E), 0x90] // U+68B5 <cjk>
	`梠`: [u8(0x9E), 0x91] // U+68A0 <cjk>
	`梺`: [u8(0x9E), 0x92] // U+68BA <cjk>
	`椏`: [u8(0x9E), 0x93] // U+690F <cjk>
	`梍`: [u8(0x9E), 0x94] // U+688D <cjk>
	`桾`: [u8(0x9E), 0x95] // U+687E <cjk>
	`椁`: [u8(0x9E), 0x96] // U+6901 <cjk>
	`棊`: [u8(0x9E), 0x97] // U+68CA <cjk>
	`椈`: [u8(0x9E), 0x98] // U+6908 <cjk>
	`棘`: [u8(0x9E), 0x99] // U+68D8 <cjk>
	`椢`: [u8(0x9E), 0x9A] // U+6922 <cjk>
	`椦`: [u8(0x9E), 0x9B] // U+6926 <cjk>
	`棡`: [u8(0x9E), 0x9C] // U+68E1 <cjk>
	`椌`: [u8(0x9E), 0x9D] // U+690C <cjk>
	`棍`: [u8(0x9E), 0x9E] // U+68CD <cjk>
	`棔`: [u8(0x9E), 0x9F] // U+68D4 <cjk>
	`棧`: [u8(0x9E), 0xA0] // U+68E7 <cjk>
	`棕`: [u8(0x9E), 0xA1] // U+68D5 <cjk>
	`椶`: [u8(0x9E), 0xA2] // U+6936 <cjk>
	`椒`: [u8(0x9E), 0xA3] // U+6912 <cjk>
	`椄`: [u8(0x9E), 0xA4] // U+6904 <cjk>
	`棗`: [u8(0x9E), 0xA5] // U+68D7 <cjk>
	`棣`: [u8(0x9E), 0xA6] // U+68E3 <cjk>
	`椥`: [u8(0x9E), 0xA7] // U+6925 <cjk>
	`棹`: [u8(0x9E), 0xA8] // U+68F9 <cjk>
	`棠`: [u8(0x9E), 0xA9] // U+68E0 <cjk>
	`棯`: [u8(0x9E), 0xAA] // U+68EF <cjk>
	`椨`: [u8(0x9E), 0xAB] // U+6928 <cjk>
	`椪`: [u8(0x9E), 0xAC] // U+692A <cjk>
	`椚`: [u8(0x9E), 0xAD] // U+691A <cjk>
	`椣`: [u8(0x9E), 0xAE] // U+6923 <cjk>
	`椡`: [u8(0x9E), 0xAF] // U+6921 <cjk>
	`棆`: [u8(0x9E), 0xB0] // U+68C6 <cjk>
	`楹`: [u8(0x9E), 0xB1] // U+6979 <cjk>
	`楷`: [u8(0x9E), 0xB2] // U+6977 <cjk>
	`楜`: [u8(0x9E), 0xB3] // U+695C <cjk>
	`楸`: [u8(0x9E), 0xB4] // U+6978 <cjk>
	`楫`: [u8(0x9E), 0xB5] // U+696B <cjk>
	`楔`: [u8(0x9E), 0xB6] // U+6954 <cjk>
	`楾`: [u8(0x9E), 0xB7] // U+697E <cjk>
	`楮`: [u8(0x9E), 0xB8] // U+696E <cjk>
	`椹`: [u8(0x9E), 0xB9] // U+6939 <cjk>
	`楴`: [u8(0x9E), 0xBA] // U+6974 <cjk>
	`椽`: [u8(0x9E), 0xBB] // U+693D <cjk>
	`楙`: [u8(0x9E), 0xBC] // U+6959 <cjk>
	`椰`: [u8(0x9E), 0xBD] // U+6930 <cjk>
	`楡`: [u8(0x9E), 0xBE] // U+6961 <cjk>
	`楞`: [u8(0x9E), 0xBF] // U+695E <cjk>
	`楝`: [u8(0x9E), 0xC0] // U+695D <cjk>
	`榁`: [u8(0x9E), 0xC1] // U+6981 <cjk>
	`楪`: [u8(0x9E), 0xC2] // U+696A <cjk>
	`榲`: [u8(0x9E), 0xC3] // U+69B2 <cjk>
	`榮`: [u8(0x9E), 0xC4] // U+69AE <cjk>
	`槐`: [u8(0x9E), 0xC5] // U+69D0 <cjk>
	`榿`: [u8(0x9E), 0xC6] // U+69BF <cjk>
	`槁`: [u8(0x9E), 0xC7] // U+69C1 <cjk>
	`槓`: [u8(0x9E), 0xC8] // U+69D3 <cjk>
	`榾`: [u8(0x9E), 0xC9] // U+69BE <cjk>
	`槎`: [u8(0x9E), 0xCA] // U+69CE <cjk>
	`寨`: [u8(0x9E), 0xCB] // U+5BE8 <cjk>
	`槊`: [u8(0x9E), 0xCC] // U+69CA <cjk>
	`槝`: [u8(0x9E), 0xCD] // U+69DD <cjk>
	`榻`: [u8(0x9E), 0xCE] // U+69BB <cjk>
	`槃`: [u8(0x9E), 0xCF] // U+69C3 <cjk>
	`榧`: [u8(0x9E), 0xD0] // U+69A7 <cjk>
	`樮`: [u8(0x9E), 0xD1] // U+6A2E <cjk>
	`榑`: [u8(0x9E), 0xD2] // U+6991 <cjk>
	`榠`: [u8(0x9E), 0xD3] // U+69A0 <cjk>
	`榜`: [u8(0x9E), 0xD4] // U+699C <cjk>
	`榕`: [u8(0x9E), 0xD5] // U+6995 <cjk>
	`榴`: [u8(0x9E), 0xD6] // U+69B4 <cjk>
	`槞`: [u8(0x9E), 0xD7] // U+69DE <cjk>
	`槨`: [u8(0x9E), 0xD8] // U+69E8 <cjk>
	`樂`: [u8(0x9E), 0xD9] // U+6A02 <cjk>
	`樛`: [u8(0x9E), 0xDA] // U+6A1B <cjk>
	`槿`: [u8(0x9E), 0xDB] // U+69FF <cjk>
	`權`: [u8(0x9E), 0xDC] // U+6B0A <cjk>
	`槹`: [u8(0x9E), 0xDD] // U+69F9 <cjk>
	`槲`: [u8(0x9E), 0xDE] // U+69F2 <cjk>
	`槧`: [u8(0x9E), 0xDF] // U+69E7 <cjk>
	`樅`: [u8(0x9E), 0xE0] // U+6A05 <cjk>
	`榱`: [u8(0x9E), 0xE1] // U+69B1 <cjk>
	`樞`: [u8(0x9E), 0xE2] // U+6A1E <cjk>
	`槭`: [u8(0x9E), 0xE3] // U+69ED <cjk>
	`樔`: [u8(0x9E), 0xE4] // U+6A14 <cjk>
	`槫`: [u8(0x9E), 0xE5] // U+69EB <cjk>
	`樊`: [u8(0x9E), 0xE6] // U+6A0A <cjk>
	`樒`: [u8(0x9E), 0xE7] // U+6A12 <cjk>
	`櫁`: [u8(0x9E), 0xE8] // U+6AC1 <cjk>
	`樣`: [u8(0x9E), 0xE9] // U+6A23 <cjk>
	`樓`: [u8(0x9E), 0xEA] // U+6A13 <cjk>
	`橄`: [u8(0x9E), 0xEB] // U+6A44 <cjk>
	`樌`: [u8(0x9E), 0xEC] // U+6A0C <cjk>
	`橲`: [u8(0x9E), 0xED] // U+6A72 <cjk>
	`樶`: [u8(0x9E), 0xEE] // U+6A36 <cjk>
	`橸`: [u8(0x9E), 0xEF] // U+6A78 <cjk>
	`橇`: [u8(0x9E), 0xF0] // U+6A47 <cjk>
	`橢`: [u8(0x9E), 0xF1] // U+6A62 <cjk>
	`橙`: [u8(0x9E), 0xF2] // U+6A59 <cjk>
	`橦`: [u8(0x9E), 0xF3] // U+6A66 <cjk>
	`橈`: [u8(0x9E), 0xF4] // U+6A48 <cjk>
	`樸`: [u8(0x9E), 0xF5] // U+6A38 <cjk>
	`樢`: [u8(0x9E), 0xF6] // U+6A22 <cjk>
	`檐`: [u8(0x9E), 0xF7] // U+6A90 <cjk>
	`檍`: [u8(0x9E), 0xF8] // U+6A8D <cjk>
	`檠`: [u8(0x9E), 0xF9] // U+6AA0 <cjk>
	`檄`: [u8(0x9E), 0xFA] // U+6A84 <cjk>
	`檢`: [u8(0x9E), 0xFB] // U+6AA2 <cjk>
	`檣`: [u8(0x9E), 0xFC] // U+6AA3 <cjk>
	`檗`: [u8(0x9F), 0x40] // U+6A97 <cjk>
	`蘗`: [u8(0x9F), 0x41] // U+8617 <cjk>
	`檻`: [u8(0x9F), 0x42] // U+6ABB <cjk>
	`櫃`: [u8(0x9F), 0x43] // U+6AC3 <cjk>
	`櫂`: [u8(0x9F), 0x44] // U+6AC2 <cjk>
	`檸`: [u8(0x9F), 0x45] // U+6AB8 <cjk>
	`檳`: [u8(0x9F), 0x46] // U+6AB3 <cjk>
	`檬`: [u8(0x9F), 0x47] // U+6AAC <cjk>
	`櫞`: [u8(0x9F), 0x48] // U+6ADE <cjk>
	`櫑`: [u8(0x9F), 0x49] // U+6AD1 <cjk>
	`櫟`: [u8(0x9F), 0x4A] // U+6ADF <cjk>
	`檪`: [u8(0x9F), 0x4B] // U+6AAA <cjk>
	`櫚`: [u8(0x9F), 0x4C] // U+6ADA <cjk>
	`櫪`: [u8(0x9F), 0x4D] // U+6AEA <cjk>
	`櫻`: [u8(0x9F), 0x4E] // U+6AFB <cjk>
	`欅`: [u8(0x9F), 0x4F] // U+6B05 <cjk>
	`蘖`: [u8(0x9F), 0x50] // U+8616 <cjk>
	`櫺`: [u8(0x9F), 0x51] // U+6AFA <cjk>
	`欒`: [u8(0x9F), 0x52] // U+6B12 <cjk>
	`欖`: [u8(0x9F), 0x53] // U+6B16 <cjk>
	`鬱`: [u8(0x9F), 0x54] // U+9B31 <cjk>
	`欟`: [u8(0x9F), 0x55] // U+6B1F <cjk>
	`欸`: [u8(0x9F), 0x56] // U+6B38 <cjk>
	`欷`: [u8(0x9F), 0x57] // U+6B37 <cjk>
	`盜`: [u8(0x9F), 0x58] // U+76DC <cjk>
	`欹`: [u8(0x9F), 0x59] // U+6B39 <cjk>
	`飮`: [u8(0x9F), 0x5A] // U+98EE <cjk>
	`歇`: [u8(0x9F), 0x5B] // U+6B47 <cjk>
	`歃`: [u8(0x9F), 0x5C] // U+6B43 <cjk>
	`歉`: [u8(0x9F), 0x5D] // U+6B49 <cjk>
	`歐`: [u8(0x9F), 0x5E] // U+6B50 <cjk>
	`歙`: [u8(0x9F), 0x5F] // U+6B59 <cjk>
	`歔`: [u8(0x9F), 0x60] // U+6B54 <cjk>
	`歛`: [u8(0x9F), 0x61] // U+6B5B <cjk>
	`歟`: [u8(0x9F), 0x62] // U+6B5F <cjk>
	`歡`: [u8(0x9F), 0x63] // U+6B61 <cjk>
	`歸`: [u8(0x9F), 0x64] // U+6B78 <cjk>
	`歹`: [u8(0x9F), 0x65] // U+6B79 <cjk>
	`歿`: [u8(0x9F), 0x66] // U+6B7F <cjk>
	`殀`: [u8(0x9F), 0x67] // U+6B80 <cjk>
	`殄`: [u8(0x9F), 0x68] // U+6B84 <cjk>
	`殃`: [u8(0x9F), 0x69] // U+6B83 <cjk>
	`殍`: [u8(0x9F), 0x6A] // U+6B8D <cjk>
	`殘`: [u8(0x9F), 0x6B] // U+6B98 <cjk>
	`殕`: [u8(0x9F), 0x6C] // U+6B95 <cjk>
	`殞`: [u8(0x9F), 0x6D] // U+6B9E <cjk>
	`殤`: [u8(0x9F), 0x6E] // U+6BA4 <cjk>
	`殪`: [u8(0x9F), 0x6F] // U+6BAA <cjk>
	`殫`: [u8(0x9F), 0x70] // U+6BAB <cjk>
	`殯`: [u8(0x9F), 0x71] // U+6BAF <cjk>
	`殲`: [u8(0x9F), 0x72] // U+6BB2 <cjk>
	`殱`: [u8(0x9F), 0x73] // U+6BB1 <cjk>
	`殳`: [u8(0x9F), 0x74] // U+6BB3 <cjk>
	`殷`: [u8(0x9F), 0x75] // U+6BB7 <cjk>
	`殼`: [u8(0x9F), 0x76] // U+6BBC <cjk>
	`毆`: [u8(0x9F), 0x77] // U+6BC6 <cjk>
	`毋`: [u8(0x9F), 0x78] // U+6BCB <cjk>
	`毓`: [u8(0x9F), 0x79] // U+6BD3 <cjk>
	`毟`: [u8(0x9F), 0x7A] // U+6BDF <cjk>
	`毬`: [u8(0x9F), 0x7B] // U+6BEC <cjk>
	`毫`: [u8(0x9F), 0x7C] // U+6BEB <cjk>
	`毳`: [u8(0x9F), 0x7D] // U+6BF3 <cjk>
	`毯`: [u8(0x9F), 0x7E] // U+6BEF <cjk>
	`麾`: [u8(0x9F), 0x80] // U+9EBE <cjk>
	`氈`: [u8(0x9F), 0x81] // U+6C08 <cjk>
	`氓`: [u8(0x9F), 0x82] // U+6C13 <cjk>
	`气`: [u8(0x9F), 0x83] // U+6C14 <cjk>
	`氛`: [u8(0x9F), 0x84] // U+6C1B <cjk>
	`氤`: [u8(0x9F), 0x85] // U+6C24 <cjk>
	`氣`: [u8(0x9F), 0x86] // U+6C23 <cjk>
	`汞`: [u8(0x9F), 0x87] // U+6C5E <cjk>
	`汕`: [u8(0x9F), 0x88] // U+6C55 <cjk>
	`汢`: [u8(0x9F), 0x89] // U+6C62 <cjk>
	`汪`: [u8(0x9F), 0x8A] // U+6C6A <cjk>
	`沂`: [u8(0x9F), 0x8B] // U+6C82 <cjk>
	`沍`: [u8(0x9F), 0x8C] // U+6C8D <cjk>
	`沚`: [u8(0x9F), 0x8D] // U+6C9A <cjk>
	`沁`: [u8(0x9F), 0x8E] // U+6C81 <cjk>
	`沛`: [u8(0x9F), 0x8F] // U+6C9B <cjk>
	`汾`: [u8(0x9F), 0x90] // U+6C7E <cjk>
	`汨`: [u8(0x9F), 0x91] // U+6C68 <cjk>
	`汳`: [u8(0x9F), 0x92] // U+6C73 <cjk>
	`沒`: [u8(0x9F), 0x93] // U+6C92 <cjk>
	`沐`: [u8(0x9F), 0x94] // U+6C90 <cjk>
	`泄`: [u8(0x9F), 0x95] // U+6CC4 <cjk>
	`泱`: [u8(0x9F), 0x96] // U+6CF1 <cjk>
	`泓`: [u8(0x9F), 0x97] // U+6CD3 <cjk>
	`沽`: [u8(0x9F), 0x98] // U+6CBD <cjk>
	`泗`: [u8(0x9F), 0x99] // U+6CD7 <cjk>
	`泅`: [u8(0x9F), 0x9A] // U+6CC5 <cjk>
	`泝`: [u8(0x9F), 0x9B] // U+6CDD <cjk>
	`沮`: [u8(0x9F), 0x9C] // U+6CAE <cjk>
	`沱`: [u8(0x9F), 0x9D] // U+6CB1 <cjk>
	`沾`: [u8(0x9F), 0x9E] // U+6CBE <cjk>
	`沺`: [u8(0x9F), 0x9F] // U+6CBA <cjk>
	`泛`: [u8(0x9F), 0xA0] // U+6CDB <cjk>
	`泯`: [u8(0x9F), 0xA1] // U+6CEF <cjk>
	`泙`: [u8(0x9F), 0xA2] // U+6CD9 <cjk>
	`泪`: [u8(0x9F), 0xA3] // U+6CEA <cjk>
	`洟`: [u8(0x9F), 0xA4] // U+6D1F <cjk>
	`衍`: [u8(0x9F), 0xA5] // U+884D <cjk>
	`洶`: [u8(0x9F), 0xA6] // U+6D36 <cjk>
	`洫`: [u8(0x9F), 0xA7] // U+6D2B <cjk>
	`洽`: [u8(0x9F), 0xA8] // U+6D3D <cjk>
	`洸`: [u8(0x9F), 0xA9] // U+6D38 <cjk>
	`洙`: [u8(0x9F), 0xAA] // U+6D19 <cjk>
	`洵`: [u8(0x9F), 0xAB] // U+6D35 <cjk>
	`洳`: [u8(0x9F), 0xAC] // U+6D33 <cjk>
	`洒`: [u8(0x9F), 0xAD] // U+6D12 <cjk>
	`洌`: [u8(0x9F), 0xAE] // U+6D0C <cjk>
	`浣`: [u8(0x9F), 0xAF] // U+6D63 <cjk>
	`涓`: [u8(0x9F), 0xB0] // U+6D93 <cjk>
	`浤`: [u8(0x9F), 0xB1] // U+6D64 <cjk>
	`浚`: [u8(0x9F), 0xB2] // U+6D5A <cjk>
	`浹`: [u8(0x9F), 0xB3] // U+6D79 <cjk>
	`浙`: [u8(0x9F), 0xB4] // U+6D59 <cjk>
	`涎`: [u8(0x9F), 0xB5] // U+6D8E <cjk>
	`涕`: [u8(0x9F), 0xB6] // U+6D95 <cjk>
	`濤`: [u8(0x9F), 0xB7] // U+6FE4 <cjk>
	`涅`: [u8(0x9F), 0xB8] // U+6D85 <cjk>
	`淹`: [u8(0x9F), 0xB9] // U+6DF9 <cjk>
	`渕`: [u8(0x9F), 0xBA] // U+6E15 <cjk>
	`渊`: [u8(0x9F), 0xBB] // U+6E0A <cjk>
	`涵`: [u8(0x9F), 0xBC] // U+6DB5 <cjk>
	`淇`: [u8(0x9F), 0xBD] // U+6DC7 <cjk>
	`淦`: [u8(0x9F), 0xBE] // U+6DE6 <cjk>
	`涸`: [u8(0x9F), 0xBF] // U+6DB8 <cjk>
	`淆`: [u8(0x9F), 0xC0] // U+6DC6 <cjk>
	`淬`: [u8(0x9F), 0xC1] // U+6DEC <cjk>
	`淞`: [u8(0x9F), 0xC2] // U+6DDE <cjk>
	`淌`: [u8(0x9F), 0xC3] // U+6DCC <cjk>
	`淨`: [u8(0x9F), 0xC4] // U+6DE8 <cjk>
	`淒`: [u8(0x9F), 0xC5] // U+6DD2 <cjk>
	`淅`: [u8(0x9F), 0xC6] // U+6DC5 <cjk>
	`淺`: [u8(0x9F), 0xC7] // U+6DFA <cjk>
	`淙`: [u8(0x9F), 0xC8] // U+6DD9 <cjk>
	`淤`: [u8(0x9F), 0xC9] // U+6DE4 <cjk>
	`淕`: [u8(0x9F), 0xCA] // U+6DD5 <cjk>
	`淪`: [u8(0x9F), 0xCB] // U+6DEA <cjk>
	`淮`: [u8(0x9F), 0xCC] // U+6DEE <cjk>
	`渭`: [u8(0x9F), 0xCD] // U+6E2D <cjk>
	`湮`: [u8(0x9F), 0xCE] // U+6E6E <cjk>
	`渮`: [u8(0x9F), 0xCF] // U+6E2E <cjk>
	`渙`: [u8(0x9F), 0xD0] // U+6E19 <cjk>
	`湲`: [u8(0x9F), 0xD1] // U+6E72 <cjk>
	`湟`: [u8(0x9F), 0xD2] // U+6E5F <cjk>
	`渾`: [u8(0x9F), 0xD3] // U+6E3E <cjk>
	`渣`: [u8(0x9F), 0xD4] // U+6E23 <cjk>
	`湫`: [u8(0x9F), 0xD5] // U+6E6B <cjk>
	`渫`: [u8(0x9F), 0xD6] // U+6E2B <cjk>
	`湶`: [u8(0x9F), 0xD7] // U+6E76 <cjk>
	`湍`: [u8(0x9F), 0xD8] // U+6E4D <cjk>
	`渟`: [u8(0x9F), 0xD9] // U+6E1F <cjk>
	`湃`: [u8(0x9F), 0xDA] // U+6E43 <cjk>
	`渺`: [u8(0x9F), 0xDB] // U+6E3A <cjk>
	`湎`: [u8(0x9F), 0xDC] // U+6E4E <cjk>
	`渤`: [u8(0x9F), 0xDD] // U+6E24 <cjk>
	`滿`: [u8(0x9F), 0xDE] // U+6EFF <cjk>
	`渝`: [u8(0x9F), 0xDF] // U+6E1D <cjk>
	`游`: [u8(0x9F), 0xE0] // U+6E38 <cjk>
	`溂`: [u8(0x9F), 0xE1] // U+6E82 <cjk>
	`溪`: [u8(0x9F), 0xE2] // U+6EAA <cjk>
	`溘`: [u8(0x9F), 0xE3] // U+6E98 <cjk>
	`滉`: [u8(0x9F), 0xE4] // U+6EC9 <cjk>
	`溷`: [u8(0x9F), 0xE5] // U+6EB7 <cjk>
	`滓`: [u8(0x9F), 0xE6] // U+6ED3 <cjk>
	`溽`: [u8(0x9F), 0xE7] // U+6EBD <cjk>
	`溯`: [u8(0x9F), 0xE8] // U+6EAF <cjk>
	`滄`: [u8(0x9F), 0xE9] // U+6EC4 <cjk>
	`溲`: [u8(0x9F), 0xEA] // U+6EB2 <cjk>
	`滔`: [u8(0x9F), 0xEB] // U+6ED4 <cjk>
	`滕`: [u8(0x9F), 0xEC] // U+6ED5 <cjk>
	`溏`: [u8(0x9F), 0xED] // U+6E8F <cjk>
	`溥`: [u8(0x9F), 0xEE] // U+6EA5 <cjk>
	`滂`: [u8(0x9F), 0xEF] // U+6EC2 <cjk>
	`溟`: [u8(0x9F), 0xF0] // U+6E9F <cjk>
	`潁`: [u8(0x9F), 0xF1] // U+6F41 <cjk>
	`漑`: [u8(0x9F), 0xF2] // U+6F11 <cjk>
	`灌`: [u8(0x9F), 0xF3] // U+704C <cjk>
	`滬`: [u8(0x9F), 0xF4] // U+6EEC <cjk>
	`滸`: [u8(0x9F), 0xF5] // U+6EF8 <cjk>
	`滾`: [u8(0x9F), 0xF6] // U+6EFE <cjk>
	`漿`: [u8(0x9F), 0xF7] // U+6F3F <cjk>
	`滲`: [u8(0x9F), 0xF8] // U+6EF2 <cjk>
	`漱`: [u8(0x9F), 0xF9] // U+6F31 <cjk>
	`滯`: [u8(0x9F), 0xFA] // U+6EEF <cjk>
	`漲`: [u8(0x9F), 0xFB] // U+6F32 <cjk>
	`滌`: [u8(0x9F), 0xFC] // U+6ECC <cjk>
	`漾`: [u8(0xE0), 0x40] // U+6F3E <cjk>
	`漓`: [u8(0xE0), 0x41] // U+6F13 <cjk>
	`滷`: [u8(0xE0), 0x42] // U+6EF7 <cjk>
	`澆`: [u8(0xE0), 0x43] // U+6F86 <cjk>
	`潺`: [u8(0xE0), 0x44] // U+6F7A <cjk>
	`潸`: [u8(0xE0), 0x45] // U+6F78 <cjk>
	`澁`: [u8(0xE0), 0x46] // U+6F81 <cjk>
	`澀`: [u8(0xE0), 0x47] // U+6F80 <cjk>
	`潯`: [u8(0xE0), 0x48] // U+6F6F <cjk>
	`潛`: [u8(0xE0), 0x49] // U+6F5B <cjk>
	`濳`: [u8(0xE0), 0x4A] // U+6FF3 <cjk>
	`潭`: [u8(0xE0), 0x4B] // U+6F6D <cjk>
	`澂`: [u8(0xE0), 0x4C] // U+6F82 <cjk>
	`潼`: [u8(0xE0), 0x4D] // U+6F7C <cjk>
	`潘`: [u8(0xE0), 0x4E] // U+6F58 <cjk>
	`澎`: [u8(0xE0), 0x4F] // U+6F8E <cjk>
	`澑`: [u8(0xE0), 0x50] // U+6F91 <cjk>
	`濂`: [u8(0xE0), 0x51] // U+6FC2 <cjk>
	`潦`: [u8(0xE0), 0x52] // U+6F66 <cjk>
	`澳`: [u8(0xE0), 0x53] // U+6FB3 <cjk>
	`澣`: [u8(0xE0), 0x54] // U+6FA3 <cjk>
	`澡`: [u8(0xE0), 0x55] // U+6FA1 <cjk>
	`澤`: [u8(0xE0), 0x56] // U+6FA4 <cjk>
	`澹`: [u8(0xE0), 0x57] // U+6FB9 <cjk>
	`濆`: [u8(0xE0), 0x58] // U+6FC6 <cjk>
	`澪`: [u8(0xE0), 0x59] // U+6FAA <cjk>
	`濟`: [u8(0xE0), 0x5A] // U+6FDF <cjk>
	`濕`: [u8(0xE0), 0x5B] // U+6FD5 <cjk>
	`濬`: [u8(0xE0), 0x5C] // U+6FEC <cjk>
	`濔`: [u8(0xE0), 0x5D] // U+6FD4 <cjk>
	`濘`: [u8(0xE0), 0x5E] // U+6FD8 <cjk>
	`濱`: [u8(0xE0), 0x5F] // U+6FF1 <cjk>
	`濮`: [u8(0xE0), 0x60] // U+6FEE <cjk>
	`濛`: [u8(0xE0), 0x61] // U+6FDB <cjk>
	`瀉`: [u8(0xE0), 0x62] // U+7009 <cjk>
	`瀋`: [u8(0xE0), 0x63] // U+700B <cjk>
	`濺`: [u8(0xE0), 0x64] // U+6FFA <cjk>
	`瀑`: [u8(0xE0), 0x65] // U+7011 <cjk>
	`瀁`: [u8(0xE0), 0x66] // U+7001 <cjk>
	`瀏`: [u8(0xE0), 0x67] // U+700F <cjk>
	`濾`: [u8(0xE0), 0x68] // U+6FFE <cjk>
	`瀛`: [u8(0xE0), 0x69] // U+701B <cjk>
	`瀚`: [u8(0xE0), 0x6A] // U+701A <cjk>
	`潴`: [u8(0xE0), 0x6B] // U+6F74 <cjk>
	`瀝`: [u8(0xE0), 0x6C] // U+701D <cjk>
	`瀘`: [u8(0xE0), 0x6D] // U+7018 <cjk>
	`瀟`: [u8(0xE0), 0x6E] // U+701F <cjk>
	`瀰`: [u8(0xE0), 0x6F] // U+7030 <cjk>
	`瀾`: [u8(0xE0), 0x70] // U+703E <cjk>
	`瀲`: [u8(0xE0), 0x71] // U+7032 <cjk>
	`灑`: [u8(0xE0), 0x72] // U+7051 <cjk>
	`灣`: [u8(0xE0), 0x73] // U+7063 <cjk>
	`炙`: [u8(0xE0), 0x74] // U+7099 <cjk>
	`炒`: [u8(0xE0), 0x75] // U+7092 <cjk>
	`炯`: [u8(0xE0), 0x76] // U+70AF <cjk>
	`烱`: [u8(0xE0), 0x77] // U+70F1 <cjk>
	`炬`: [u8(0xE0), 0x78] // U+70AC <cjk>
	`炸`: [u8(0xE0), 0x79] // U+70B8 <cjk>
	`炳`: [u8(0xE0), 0x7A] // U+70B3 <cjk>
	`炮`: [u8(0xE0), 0x7B] // U+70AE <cjk>
	`烟`: [u8(0xE0), 0x7C] // U+70DF <cjk>
	`烋`: [u8(0xE0), 0x7D] // U+70CB <cjk>
	`烝`: [u8(0xE0), 0x7E] // U+70DD <cjk>
	`烙`: [u8(0xE0), 0x80] // U+70D9 <cjk>
	`焉`: [u8(0xE0), 0x81] // U+7109 <cjk>
	`烽`: [u8(0xE0), 0x82] // U+70FD <cjk>
	`焜`: [u8(0xE0), 0x83] // U+711C <cjk>
	`焙`: [u8(0xE0), 0x84] // U+7119 <cjk>
	`煥`: [u8(0xE0), 0x85] // U+7165 <cjk>
	`煕`: [u8(0xE0), 0x86] // U+7155 <cjk>
	`熈`: [u8(0xE0), 0x87] // U+7188 <cjk>
	`煦`: [u8(0xE0), 0x88] // U+7166 <cjk>
	`煢`: [u8(0xE0), 0x89] // U+7162 <cjk>
	`煌`: [u8(0xE0), 0x8A] // U+714C <cjk>
	`煖`: [u8(0xE0), 0x8B] // U+7156 <cjk>
	`煬`: [u8(0xE0), 0x8C] // U+716C <cjk>
	`熏`: [u8(0xE0), 0x8D] // U+718F <cjk>
	`燻`: [u8(0xE0), 0x8E] // U+71FB <cjk>
	`熄`: [u8(0xE0), 0x8F] // U+7184 <cjk>
	`熕`: [u8(0xE0), 0x90] // U+7195 <cjk>
	`熨`: [u8(0xE0), 0x91] // U+71A8 <cjk>
	`熬`: [u8(0xE0), 0x92] // U+71AC <cjk>
	`燗`: [u8(0xE0), 0x93] // U+71D7 <cjk>
	`熹`: [u8(0xE0), 0x94] // U+71B9 <cjk>
	`熾`: [u8(0xE0), 0x95] // U+71BE <cjk>
	`燒`: [u8(0xE0), 0x96] // U+71D2 <cjk>
	`燉`: [u8(0xE0), 0x97] // U+71C9 <cjk>
	`燔`: [u8(0xE0), 0x98] // U+71D4 <cjk>
	`燎`: [u8(0xE0), 0x99] // U+71CE <cjk>
	`燠`: [u8(0xE0), 0x9A] // U+71E0 <cjk>
	`燬`: [u8(0xE0), 0x9B] // U+71EC <cjk>
	`燧`: [u8(0xE0), 0x9C] // U+71E7 <cjk>
	`燵`: [u8(0xE0), 0x9D] // U+71F5 <cjk>
	`燼`: [u8(0xE0), 0x9E] // U+71FC <cjk>
	`燹`: [u8(0xE0), 0x9F] // U+71F9 <cjk>
	`燿`: [u8(0xE0), 0xA0] // U+71FF <cjk>
	`爍`: [u8(0xE0), 0xA1] // U+720D <cjk>
	`爐`: [u8(0xE0), 0xA2] // U+7210 <cjk>
	`爛`: [u8(0xE0), 0xA3] // U+721B <cjk>
	`爨`: [u8(0xE0), 0xA4] // U+7228 <cjk>
	`爭`: [u8(0xE0), 0xA5] // U+722D <cjk>
	`爬`: [u8(0xE0), 0xA6] // U+722C <cjk>
	`爰`: [u8(0xE0), 0xA7] // U+7230 <cjk>
	`爲`: [u8(0xE0), 0xA8] // U+7232 <cjk>
	`爻`: [u8(0xE0), 0xA9] // U+723B <cjk>
	`爼`: [u8(0xE0), 0xAA] // U+723C <cjk>
	`爿`: [u8(0xE0), 0xAB] // U+723F <cjk>
	`牀`: [u8(0xE0), 0xAC] // U+7240 <cjk>
	`牆`: [u8(0xE0), 0xAD] // U+7246 <cjk>
	`牋`: [u8(0xE0), 0xAE] // U+724B <cjk>
	`牘`: [u8(0xE0), 0xAF] // U+7258 <cjk>
	`牴`: [u8(0xE0), 0xB0] // U+7274 <cjk>
	`牾`: [u8(0xE0), 0xB1] // U+727E <cjk>
	`犂`: [u8(0xE0), 0xB2] // U+7282 <cjk>
	`犁`: [u8(0xE0), 0xB3] // U+7281 <cjk>
	`犇`: [u8(0xE0), 0xB4] // U+7287 <cjk>
	`犒`: [u8(0xE0), 0xB5] // U+7292 <cjk>
	`犖`: [u8(0xE0), 0xB6] // U+7296 <cjk>
	`犢`: [u8(0xE0), 0xB7] // U+72A2 <cjk>
	`犧`: [u8(0xE0), 0xB8] // U+72A7 <cjk>
	`犹`: [u8(0xE0), 0xB9] // U+72B9 <cjk>
	`犲`: [u8(0xE0), 0xBA] // U+72B2 <cjk>
	`狃`: [u8(0xE0), 0xBB] // U+72C3 <cjk>
	`狆`: [u8(0xE0), 0xBC] // U+72C6 <cjk>
	`狄`: [u8(0xE0), 0xBD] // U+72C4 <cjk>
	`狎`: [u8(0xE0), 0xBE] // U+72CE <cjk>
	`狒`: [u8(0xE0), 0xBF] // U+72D2 <cjk>
	`狢`: [u8(0xE0), 0xC0] // U+72E2 <cjk>
	`狠`: [u8(0xE0), 0xC1] // U+72E0 <cjk>
	`狡`: [u8(0xE0), 0xC2] // U+72E1 <cjk>
	`狹`: [u8(0xE0), 0xC3] // U+72F9 <cjk>
	`狷`: [u8(0xE0), 0xC4] // U+72F7 <cjk>
	`倏`: [u8(0xE0), 0xC5] // U+500F <cjk>
	`猗`: [u8(0xE0), 0xC6] // U+7317 <cjk>
	`猊`: [u8(0xE0), 0xC7] // U+730A <cjk>
	`猜`: [u8(0xE0), 0xC8] // U+731C <cjk>
	`猖`: [u8(0xE0), 0xC9] // U+7316 <cjk>
	`猝`: [u8(0xE0), 0xCA] // U+731D <cjk>
	`猴`: [u8(0xE0), 0xCB] // U+7334 <cjk>
	`猯`: [u8(0xE0), 0xCC] // U+732F <cjk>
	`猩`: [u8(0xE0), 0xCD] // U+7329 <cjk>
	`猥`: [u8(0xE0), 0xCE] // U+7325 <cjk>
	`猾`: [u8(0xE0), 0xCF] // U+733E <cjk>
	`獎`: [u8(0xE0), 0xD0] // U+734E <cjk>
	`獏`: [u8(0xE0), 0xD1] // U+734F <cjk>
	`默`: [u8(0xE0), 0xD2] // U+9ED8 <cjk>
	`獗`: [u8(0xE0), 0xD3] // U+7357 <cjk>
	`獪`: [u8(0xE0), 0xD4] // U+736A <cjk>
	`獨`: [u8(0xE0), 0xD5] // U+7368 <cjk>
	`獰`: [u8(0xE0), 0xD6] // U+7370 <cjk>
	`獸`: [u8(0xE0), 0xD7] // U+7378 <cjk>
	`獵`: [u8(0xE0), 0xD8] // U+7375 <cjk>
	`獻`: [u8(0xE0), 0xD9] // U+737B <cjk>
	`獺`: [u8(0xE0), 0xDA] // U+737A <cjk>
	`珈`: [u8(0xE0), 0xDB] // U+73C8 <cjk>
	`玳`: [u8(0xE0), 0xDC] // U+73B3 <cjk>
	`珎`: [u8(0xE0), 0xDD] // U+73CE <cjk>
	`玻`: [u8(0xE0), 0xDE] // U+73BB <cjk>
	`珀`: [u8(0xE0), 0xDF] // U+73C0 <cjk>
	`珥`: [u8(0xE0), 0xE0] // U+73E5 <cjk>
	`珮`: [u8(0xE0), 0xE1] // U+73EE <cjk>
	`珞`: [u8(0xE0), 0xE2] // U+73DE <cjk>
	`璢`: [u8(0xE0), 0xE3] // U+74A2 <cjk>
	`琅`: [u8(0xE0), 0xE4] // U+7405 <cjk>
	`瑯`: [u8(0xE0), 0xE5] // U+746F <cjk>
	`琥`: [u8(0xE0), 0xE6] // U+7425 <cjk>
	`珸`: [u8(0xE0), 0xE7] // U+73F8 <cjk>
	`琲`: [u8(0xE0), 0xE8] // U+7432 <cjk>
	`琺`: [u8(0xE0), 0xE9] // U+743A <cjk>
	`瑕`: [u8(0xE0), 0xEA] // U+7455 <cjk>
	`琿`: [u8(0xE0), 0xEB] // U+743F <cjk>
	`瑟`: [u8(0xE0), 0xEC] // U+745F <cjk>
	`瑙`: [u8(0xE0), 0xED] // U+7459 <cjk>
	`瑁`: [u8(0xE0), 0xEE] // U+7441 <cjk>
	`瑜`: [u8(0xE0), 0xEF] // U+745C <cjk>
	`瑩`: [u8(0xE0), 0xF0] // U+7469 <cjk>
	`瑰`: [u8(0xE0), 0xF1] // U+7470 <cjk>
	`瑣`: [u8(0xE0), 0xF2] // U+7463 <cjk>
	`瑪`: [u8(0xE0), 0xF3] // U+746A <cjk>
	`瑶`: [u8(0xE0), 0xF4] // U+7476 <cjk>
	`瑾`: [u8(0xE0), 0xF5] // U+747E <cjk>
	`璋`: [u8(0xE0), 0xF6] // U+748B <cjk>
	`璞`: [u8(0xE0), 0xF7] // U+749E <cjk>
	`璧`: [u8(0xE0), 0xF8] // U+74A7 <cjk>
	`瓊`: [u8(0xE0), 0xF9] // U+74CA <cjk>
	`瓏`: [u8(0xE0), 0xFA] // U+74CF <cjk>
	`瓔`: [u8(0xE0), 0xFB] // U+74D4 <cjk>
	`珱`: [u8(0xE0), 0xFC] // U+73F1 <cjk>
	`瓠`: [u8(0xE1), 0x40] // U+74E0 <cjk>
	`瓣`: [u8(0xE1), 0x41] // U+74E3 <cjk>
	`瓧`: [u8(0xE1), 0x42] // U+74E7 <cjk>
	`瓩`: [u8(0xE1), 0x43] // U+74E9 <cjk>
	`瓮`: [u8(0xE1), 0x44] // U+74EE <cjk>
	`瓲`: [u8(0xE1), 0x45] // U+74F2 <cjk>
	`瓰`: [u8(0xE1), 0x46] // U+74F0 <cjk>
	`瓱`: [u8(0xE1), 0x47] // U+74F1 <cjk>
	`瓸`: [u8(0xE1), 0x48] // U+74F8 <cjk>
	`瓷`: [u8(0xE1), 0x49] // U+74F7 <cjk>
	`甄`: [u8(0xE1), 0x4A] // U+7504 <cjk>
	`甃`: [u8(0xE1), 0x4B] // U+7503 <cjk>
	`甅`: [u8(0xE1), 0x4C] // U+7505 <cjk>
	`甌`: [u8(0xE1), 0x4D] // U+750C <cjk>
	`甎`: [u8(0xE1), 0x4E] // U+750E <cjk>
	`甍`: [u8(0xE1), 0x4F] // U+750D <cjk>
	`甕`: [u8(0xE1), 0x50] // U+7515 <cjk>
	`甓`: [u8(0xE1), 0x51] // U+7513 <cjk>
	`甞`: [u8(0xE1), 0x52] // U+751E <cjk>
	`甦`: [u8(0xE1), 0x53] // U+7526 <cjk>
	`甬`: [u8(0xE1), 0x54] // U+752C <cjk>
	`甼`: [u8(0xE1), 0x55] // U+753C <cjk>
	`畄`: [u8(0xE1), 0x56] // U+7544 <cjk>
	`畍`: [u8(0xE1), 0x57] // U+754D <cjk>
	`畊`: [u8(0xE1), 0x58] // U+754A <cjk>
	`畉`: [u8(0xE1), 0x59] // U+7549 <cjk>
	`畛`: [u8(0xE1), 0x5A] // U+755B <cjk>
	`畆`: [u8(0xE1), 0x5B] // U+7546 <cjk>
	`畚`: [u8(0xE1), 0x5C] // U+755A <cjk>
	`畩`: [u8(0xE1), 0x5D] // U+7569 <cjk>
	`畤`: [u8(0xE1), 0x5E] // U+7564 <cjk>
	`畧`: [u8(0xE1), 0x5F] // U+7567 <cjk>
	`畫`: [u8(0xE1), 0x60] // U+756B <cjk>
	`畭`: [u8(0xE1), 0x61] // U+756D <cjk>
	`畸`: [u8(0xE1), 0x62] // U+7578 <cjk>
	`當`: [u8(0xE1), 0x63] // U+7576 <cjk>
	`疆`: [u8(0xE1), 0x64] // U+7586 <cjk>
	`疇`: [u8(0xE1), 0x65] // U+7587 <cjk>
	`畴`: [u8(0xE1), 0x66] // U+7574 <cjk>
	`疊`: [u8(0xE1), 0x67] // U+758A <cjk>
	`疉`: [u8(0xE1), 0x68] // U+7589 <cjk>
	`疂`: [u8(0xE1), 0x69] // U+7582 <cjk>
	`疔`: [u8(0xE1), 0x6A] // U+7594 <cjk>
	`疚`: [u8(0xE1), 0x6B] // U+759A <cjk>
	`疝`: [u8(0xE1), 0x6C] // U+759D <cjk>
	`疥`: [u8(0xE1), 0x6D] // U+75A5 <cjk>
	`疣`: [u8(0xE1), 0x6E] // U+75A3 <cjk>
	`痂`: [u8(0xE1), 0x6F] // U+75C2 <cjk>
	`疳`: [u8(0xE1), 0x70] // U+75B3 <cjk>
	`痃`: [u8(0xE1), 0x71] // U+75C3 <cjk>
	`疵`: [u8(0xE1), 0x72] // U+75B5 <cjk>
	`疽`: [u8(0xE1), 0x73] // U+75BD <cjk>
	`疸`: [u8(0xE1), 0x74] // U+75B8 <cjk>
	`疼`: [u8(0xE1), 0x75] // U+75BC <cjk>
	`疱`: [u8(0xE1), 0x76] // U+75B1 <cjk>
	`痍`: [u8(0xE1), 0x77] // U+75CD <cjk>
	`痊`: [u8(0xE1), 0x78] // U+75CA <cjk>
	`痒`: [u8(0xE1), 0x79] // U+75D2 <cjk>
	`痙`: [u8(0xE1), 0x7A] // U+75D9 <cjk>
	`痣`: [u8(0xE1), 0x7B] // U+75E3 <cjk>
	`痞`: [u8(0xE1), 0x7C] // U+75DE <cjk>
	`痾`: [u8(0xE1), 0x7D] // U+75FE <cjk>
	`痿`: [u8(0xE1), 0x7E] // U+75FF <cjk>
	`痼`: [u8(0xE1), 0x80] // U+75FC <cjk>
	`瘁`: [u8(0xE1), 0x81] // U+7601 <cjk>
	`痰`: [u8(0xE1), 0x82] // U+75F0 <cjk>
	`痺`: [u8(0xE1), 0x83] // U+75FA <cjk>
	`痲`: [u8(0xE1), 0x84] // U+75F2 <cjk>
	`痳`: [u8(0xE1), 0x85] // U+75F3 <cjk>
	`瘋`: [u8(0xE1), 0x86] // U+760B <cjk>
	`瘍`: [u8(0xE1), 0x87] // U+760D <cjk>
	`瘉`: [u8(0xE1), 0x88] // U+7609 <cjk>
	`瘟`: [u8(0xE1), 0x89] // U+761F <cjk>
	`瘧`: [u8(0xE1), 0x8A] // U+7627 <cjk>
	`瘠`: [u8(0xE1), 0x8B] // U+7620 <cjk>
	`瘡`: [u8(0xE1), 0x8C] // U+7621 <cjk>
	`瘢`: [u8(0xE1), 0x8D] // U+7622 <cjk>
	`瘤`: [u8(0xE1), 0x8E] // U+7624 <cjk>
	`瘴`: [u8(0xE1), 0x8F] // U+7634 <cjk>
	`瘰`: [u8(0xE1), 0x90] // U+7630 <cjk>
	`瘻`: [u8(0xE1), 0x91] // U+763B <cjk>
	`癇`: [u8(0xE1), 0x92] // U+7647 <cjk>
	`癈`: [u8(0xE1), 0x93] // U+7648 <cjk>
	`癆`: [u8(0xE1), 0x94] // U+7646 <cjk>
	`癜`: [u8(0xE1), 0x95] // U+765C <cjk>
	`癘`: [u8(0xE1), 0x96] // U+7658 <cjk>
	`癡`: [u8(0xE1), 0x97] // U+7661 <cjk>
	`癢`: [u8(0xE1), 0x98] // U+7662 <cjk>
	`癨`: [u8(0xE1), 0x99] // U+7668 <cjk>
	`癩`: [u8(0xE1), 0x9A] // U+7669 <cjk>
	`癪`: [u8(0xE1), 0x9B] // U+766A <cjk>
	`癧`: [u8(0xE1), 0x9C] // U+7667 <cjk>
	`癬`: [u8(0xE1), 0x9D] // U+766C <cjk>
	`癰`: [u8(0xE1), 0x9E] // U+7670 <cjk>
	`癲`: [u8(0xE1), 0x9F] // U+7672 <cjk>
	`癶`: [u8(0xE1), 0xA0] // U+7676 <cjk>
	`癸`: [u8(0xE1), 0xA1] // U+7678 <cjk>
	`發`: [u8(0xE1), 0xA2] // U+767C <cjk>
	`皀`: [u8(0xE1), 0xA3] // U+7680 <cjk>
	`皃`: [u8(0xE1), 0xA4] // U+7683 <cjk>
	`皈`: [u8(0xE1), 0xA5] // U+7688 <cjk>
	`皋`: [u8(0xE1), 0xA6] // U+768B <cjk>
	`皎`: [u8(0xE1), 0xA7] // U+768E <cjk>
	`皖`: [u8(0xE1), 0xA8] // U+7696 <cjk>
	`皓`: [u8(0xE1), 0xA9] // U+7693 <cjk>
	`皙`: [u8(0xE1), 0xAA] // U+7699 <cjk>
	`皚`: [u8(0xE1), 0xAB] // U+769A <cjk>
	`皰`: [u8(0xE1), 0xAC] // U+76B0 <cjk>
	`皴`: [u8(0xE1), 0xAD] // U+76B4 <cjk>
	`皸`: [u8(0xE1), 0xAE] // U+76B8 <cjk>
	`皹`: [u8(0xE1), 0xAF] // U+76B9 <cjk>
	`皺`: [u8(0xE1), 0xB0] // U+76BA <cjk>
	`盂`: [u8(0xE1), 0xB1] // U+76C2 <cjk>
	`盍`: [u8(0xE1), 0xB2] // U+76CD <cjk>
	`盖`: [u8(0xE1), 0xB3] // U+76D6 <cjk>
	`盒`: [u8(0xE1), 0xB4] // U+76D2 <cjk>
	`盞`: [u8(0xE1), 0xB5] // U+76DE <cjk>
	`盡`: [u8(0xE1), 0xB6] // U+76E1 <cjk>
	`盥`: [u8(0xE1), 0xB7] // U+76E5 <cjk>
	`盧`: [u8(0xE1), 0xB8] // U+76E7 <cjk>
	`盪`: [u8(0xE1), 0xB9] // U+76EA <cjk>
	`蘯`: [u8(0xE1), 0xBA] // U+862F <cjk>
	`盻`: [u8(0xE1), 0xBB] // U+76FB <cjk>
	`眈`: [u8(0xE1), 0xBC] // U+7708 <cjk>
	`眇`: [u8(0xE1), 0xBD] // U+7707 <cjk>
	`眄`: [u8(0xE1), 0xBE] // U+7704 <cjk>
	`眩`: [u8(0xE1), 0xBF] // U+7729 <cjk>
	`眤`: [u8(0xE1), 0xC0] // U+7724 <cjk>
	`眞`: [u8(0xE1), 0xC1] // U+771E <cjk>
	`眥`: [u8(0xE1), 0xC2] // U+7725 <cjk>
	`眦`: [u8(0xE1), 0xC3] // U+7726 <cjk>
	`眛`: [u8(0xE1), 0xC4] // U+771B <cjk>
	`眷`: [u8(0xE1), 0xC5] // U+7737 <cjk>
	`眸`: [u8(0xE1), 0xC6] // U+7738 <cjk>
	`睇`: [u8(0xE1), 0xC7] // U+7747 <cjk>
	`睚`: [u8(0xE1), 0xC8] // U+775A <cjk>
	`睨`: [u8(0xE1), 0xC9] // U+7768 <cjk>
	`睫`: [u8(0xE1), 0xCA] // U+776B <cjk>
	`睛`: [u8(0xE1), 0xCB] // U+775B <cjk>
	`睥`: [u8(0xE1), 0xCC] // U+7765 <cjk>
	`睿`: [u8(0xE1), 0xCD] // U+777F <cjk>
	`睾`: [u8(0xE1), 0xCE] // U+777E <cjk>
	`睹`: [u8(0xE1), 0xCF] // U+7779 <cjk>
	`瞎`: [u8(0xE1), 0xD0] // U+778E <cjk>
	`瞋`: [u8(0xE1), 0xD1] // U+778B <cjk>
	`瞑`: [u8(0xE1), 0xD2] // U+7791 <cjk>
	`瞠`: [u8(0xE1), 0xD3] // U+77A0 <cjk>
	`瞞`: [u8(0xE1), 0xD4] // U+779E <cjk>
	`瞰`: [u8(0xE1), 0xD5] // U+77B0 <cjk>
	`瞶`: [u8(0xE1), 0xD6] // U+77B6 <cjk>
	`瞹`: [u8(0xE1), 0xD7] // U+77B9 <cjk>
	`瞿`: [u8(0xE1), 0xD8] // U+77BF <cjk>
	`瞼`: [u8(0xE1), 0xD9] // U+77BC <cjk>
	`瞽`: [u8(0xE1), 0xDA] // U+77BD <cjk>
	`瞻`: [u8(0xE1), 0xDB] // U+77BB <cjk>
	`矇`: [u8(0xE1), 0xDC] // U+77C7 <cjk>
	`矍`: [u8(0xE1), 0xDD] // U+77CD <cjk>
	`矗`: [u8(0xE1), 0xDE] // U+77D7 <cjk>
	`矚`: [u8(0xE1), 0xDF] // U+77DA <cjk>
	`矜`: [u8(0xE1), 0xE0] // U+77DC <cjk>
	`矣`: [u8(0xE1), 0xE1] // U+77E3 <cjk>
	`矮`: [u8(0xE1), 0xE2] // U+77EE <cjk>
	`矼`: [u8(0xE1), 0xE3] // U+77FC <cjk>
	`砌`: [u8(0xE1), 0xE4] // U+780C <cjk>
	`砒`: [u8(0xE1), 0xE5] // U+7812 <cjk>
	`礦`: [u8(0xE1), 0xE6] // U+7926 <cjk>
	`砠`: [u8(0xE1), 0xE7] // U+7820 <cjk>
	`礪`: [u8(0xE1), 0xE8] // U+792A <cjk>
	`硅`: [u8(0xE1), 0xE9] // U+7845 <cjk>
	`碎`: [u8(0xE1), 0xEA] // U+788E <cjk>
	`硴`: [u8(0xE1), 0xEB] // U+7874 <cjk>
	`碆`: [u8(0xE1), 0xEC] // U+7886 <cjk>
	`硼`: [u8(0xE1), 0xED] // U+787C <cjk>
	`碚`: [u8(0xE1), 0xEE] // U+789A <cjk>
	`碌`: [u8(0xE1), 0xEF] // U+788C <cjk>
	`碣`: [u8(0xE1), 0xF0] // U+78A3 <cjk>
	`碵`: [u8(0xE1), 0xF1] // U+78B5 <cjk>
	`碪`: [u8(0xE1), 0xF2] // U+78AA <cjk>
	`碯`: [u8(0xE1), 0xF3] // U+78AF <cjk>
	`磑`: [u8(0xE1), 0xF4] // U+78D1 <cjk>
	`磆`: [u8(0xE1), 0xF5] // U+78C6 <cjk>
	`磋`: [u8(0xE1), 0xF6] // U+78CB <cjk>
	`磔`: [u8(0xE1), 0xF7] // U+78D4 <cjk>
	`碾`: [u8(0xE1), 0xF8] // U+78BE <cjk>
	`碼`: [u8(0xE1), 0xF9] // U+78BC <cjk>
	`磅`: [u8(0xE1), 0xFA] // U+78C5 <cjk>
	`磊`: [u8(0xE1), 0xFB] // U+78CA <cjk>
	`磬`: [u8(0xE1), 0xFC] // U+78EC <cjk>
	`磧`: [u8(0xE2), 0x40] // U+78E7 <cjk>
	`磚`: [u8(0xE2), 0x41] // U+78DA <cjk>
	`磽`: [u8(0xE2), 0x42] // U+78FD <cjk>
	`磴`: [u8(0xE2), 0x43] // U+78F4 <cjk>
	`礇`: [u8(0xE2), 0x44] // U+7907 <cjk>
	`礒`: [u8(0xE2), 0x45] // U+7912 <cjk>
	`礑`: [u8(0xE2), 0x46] // U+7911 <cjk>
	`礙`: [u8(0xE2), 0x47] // U+7919 <cjk>
	`礬`: [u8(0xE2), 0x48] // U+792C <cjk>
	`礫`: [u8(0xE2), 0x49] // U+792B <cjk>
	`祀`: [u8(0xE2), 0x4A] // U+7940 <cjk>
	`祠`: [u8(0xE2), 0x4B] // U+7960 <cjk>
	`祗`: [u8(0xE2), 0x4C] // U+7957 <cjk>
	`祟`: [u8(0xE2), 0x4D] // U+795F <cjk>
	`祚`: [u8(0xE2), 0x4E] // U+795A <cjk>
	`祕`: [u8(0xE2), 0x4F] // U+7955 <cjk>
	`祓`: [u8(0xE2), 0x50] // U+7953 <cjk>
	`祺`: [u8(0xE2), 0x51] // U+797A <cjk>
	`祿`: [u8(0xE2), 0x52] // U+797F <cjk>
	`禊`: [u8(0xE2), 0x53] // U+798A <cjk>
	`禝`: [u8(0xE2), 0x54] // U+799D <cjk>
	`禧`: [u8(0xE2), 0x55] // U+79A7 <cjk>
	`齋`: [u8(0xE2), 0x56] // U+9F4B <cjk>
	`禪`: [u8(0xE2), 0x57] // U+79AA <cjk>
	`禮`: [u8(0xE2), 0x58] // U+79AE <cjk>
	`禳`: [u8(0xE2), 0x59] // U+79B3 <cjk>
	`禹`: [u8(0xE2), 0x5A] // U+79B9 <cjk>
	`禺`: [u8(0xE2), 0x5B] // U+79BA <cjk>
	`秉`: [u8(0xE2), 0x5C] // U+79C9 <cjk>
	`秕`: [u8(0xE2), 0x5D] // U+79D5 <cjk>
	`秧`: [u8(0xE2), 0x5E] // U+79E7 <cjk>
	`秬`: [u8(0xE2), 0x5F] // U+79EC <cjk>
	`秡`: [u8(0xE2), 0x60] // U+79E1 <cjk>
	`秣`: [u8(0xE2), 0x61] // U+79E3 <cjk>
	`稈`: [u8(0xE2), 0x62] // U+7A08 <cjk>
	`稍`: [u8(0xE2), 0x63] // U+7A0D <cjk>
	`稘`: [u8(0xE2), 0x64] // U+7A18 <cjk>
	`稙`: [u8(0xE2), 0x65] // U+7A19 <cjk>
	`稠`: [u8(0xE2), 0x66] // U+7A20 <cjk>
	`稟`: [u8(0xE2), 0x67] // U+7A1F <cjk>
	`禀`: [u8(0xE2), 0x68] // U+7980 <cjk>
	`稱`: [u8(0xE2), 0x69] // U+7A31 <cjk>
	`稻`: [u8(0xE2), 0x6A] // U+7A3B <cjk>
	`稾`: [u8(0xE2), 0x6B] // U+7A3E <cjk>
	`稷`: [u8(0xE2), 0x6C] // U+7A37 <cjk>
	`穃`: [u8(0xE2), 0x6D] // U+7A43 <cjk>
	`穗`: [u8(0xE2), 0x6E] // U+7A57 <cjk>
	`穉`: [u8(0xE2), 0x6F] // U+7A49 <cjk>
	`穡`: [u8(0xE2), 0x70] // U+7A61 <cjk>
	`穢`: [u8(0xE2), 0x71] // U+7A62 <cjk>
	`穩`: [u8(0xE2), 0x72] // U+7A69 <cjk>
	`龝`: [u8(0xE2), 0x73] // U+9F9D <cjk>
	`穰`: [u8(0xE2), 0x74] // U+7A70 <cjk>
	`穹`: [u8(0xE2), 0x75] // U+7A79 <cjk>
	`穽`: [u8(0xE2), 0x76] // U+7A7D <cjk>
	`窈`: [u8(0xE2), 0x77] // U+7A88 <cjk>
	`窗`: [u8(0xE2), 0x78] // U+7A97 <cjk>
	`窕`: [u8(0xE2), 0x79] // U+7A95 <cjk>
	`窘`: [u8(0xE2), 0x7A] // U+7A98 <cjk>
	`窖`: [u8(0xE2), 0x7B] // U+7A96 <cjk>
	`窩`: [u8(0xE2), 0x7C] // U+7AA9 <cjk>
	`竈`: [u8(0xE2), 0x7D] // U+7AC8 <cjk>
	`窰`: [u8(0xE2), 0x7E] // U+7AB0 <cjk>
	`窶`: [u8(0xE2), 0x80] // U+7AB6 <cjk>
	`竅`: [u8(0xE2), 0x81] // U+7AC5 <cjk>
	`竄`: [u8(0xE2), 0x82] // U+7AC4 <cjk>
	`窿`: [u8(0xE2), 0x83] // U+7ABF <cjk>
	`邃`: [u8(0xE2), 0x84] // U+9083 <cjk>
	`竇`: [u8(0xE2), 0x85] // U+7AC7 <cjk>
	`竊`: [u8(0xE2), 0x86] // U+7ACA <cjk>
	`竍`: [u8(0xE2), 0x87] // U+7ACD <cjk>
	`竏`: [u8(0xE2), 0x88] // U+7ACF <cjk>
	`竕`: [u8(0xE2), 0x89] // U+7AD5 <cjk>
	`竓`: [u8(0xE2), 0x8A] // U+7AD3 <cjk>
	`站`: [u8(0xE2), 0x8B] // U+7AD9 <cjk>
	`竚`: [u8(0xE2), 0x8C] // U+7ADA <cjk>
	`竝`: [u8(0xE2), 0x8D] // U+7ADD <cjk>
	`竡`: [u8(0xE2), 0x8E] // U+7AE1 <cjk>
	`竢`: [u8(0xE2), 0x8F] // U+7AE2 <cjk>
	`竦`: [u8(0xE2), 0x90] // U+7AE6 <cjk>
	`竭`: [u8(0xE2), 0x91] // U+7AED <cjk>
	`竰`: [u8(0xE2), 0x92] // U+7AF0 <cjk>
	`笂`: [u8(0xE2), 0x93] // U+7B02 <cjk>
	`笏`: [u8(0xE2), 0x94] // U+7B0F <cjk>
	`笊`: [u8(0xE2), 0x95] // U+7B0A <cjk>
	`笆`: [u8(0xE2), 0x96] // U+7B06 <cjk>
	`笳`: [u8(0xE2), 0x97] // U+7B33 <cjk>
	`笘`: [u8(0xE2), 0x98] // U+7B18 <cjk>
	`笙`: [u8(0xE2), 0x99] // U+7B19 <cjk>
	`笞`: [u8(0xE2), 0x9A] // U+7B1E <cjk>
	`笵`: [u8(0xE2), 0x9B] // U+7B35 <cjk>
	`笨`: [u8(0xE2), 0x9C] // U+7B28 <cjk>
	`笶`: [u8(0xE2), 0x9D] // U+7B36 <cjk>
	`筐`: [u8(0xE2), 0x9E] // U+7B50 <cjk>
	`筺`: [u8(0xE2), 0x9F] // U+7B7A <cjk>
	`笄`: [u8(0xE2), 0xA0] // U+7B04 <cjk>
	`筍`: [u8(0xE2), 0xA1] // U+7B4D <cjk>
	`笋`: [u8(0xE2), 0xA2] // U+7B0B <cjk>
	`筌`: [u8(0xE2), 0xA3] // U+7B4C <cjk>
	`筅`: [u8(0xE2), 0xA4] // U+7B45 <cjk>
	`筵`: [u8(0xE2), 0xA5] // U+7B75 <cjk>
	`筥`: [u8(0xE2), 0xA6] // U+7B65 <cjk>
	`筴`: [u8(0xE2), 0xA7] // U+7B74 <cjk>
	`筧`: [u8(0xE2), 0xA8] // U+7B67 <cjk>
	`筰`: [u8(0xE2), 0xA9] // U+7B70 <cjk>
	`筱`: [u8(0xE2), 0xAA] // U+7B71 <cjk>
	`筬`: [u8(0xE2), 0xAB] // U+7B6C <cjk>
	`筮`: [u8(0xE2), 0xAC] // U+7B6E <cjk>
	`箝`: [u8(0xE2), 0xAD] // U+7B9D <cjk>
	`箘`: [u8(0xE2), 0xAE] // U+7B98 <cjk>
	`箟`: [u8(0xE2), 0xAF] // U+7B9F <cjk>
	`箍`: [u8(0xE2), 0xB0] // U+7B8D <cjk>
	`箜`: [u8(0xE2), 0xB1] // U+7B9C <cjk>
	`箚`: [u8(0xE2), 0xB2] // U+7B9A <cjk>
	`箋`: [u8(0xE2), 0xB3] // U+7B8B <cjk>
	`箒`: [u8(0xE2), 0xB4] // U+7B92 <cjk>
	`箏`: [u8(0xE2), 0xB5] // U+7B8F <cjk>
	`筝`: [u8(0xE2), 0xB6] // U+7B5D <cjk>
	`箙`: [u8(0xE2), 0xB7] // U+7B99 <cjk>
	`篋`: [u8(0xE2), 0xB8] // U+7BCB <cjk>
	`篁`: [u8(0xE2), 0xB9] // U+7BC1 <cjk>
	`篌`: [u8(0xE2), 0xBA] // U+7BCC <cjk>
	`篏`: [u8(0xE2), 0xBB] // U+7BCF <cjk>
	`箴`: [u8(0xE2), 0xBC] // U+7BB4 <cjk>
	`篆`: [u8(0xE2), 0xBD] // U+7BC6 <cjk>
	`篝`: [u8(0xE2), 0xBE] // U+7BDD <cjk>
	`篩`: [u8(0xE2), 0xBF] // U+7BE9 <cjk>
	`簑`: [u8(0xE2), 0xC0] // U+7C11 <cjk>
	`簔`: [u8(0xE2), 0xC1] // U+7C14 <cjk>
	`篦`: [u8(0xE2), 0xC2] // U+7BE6 <cjk>
	`篥`: [u8(0xE2), 0xC3] // U+7BE5 <cjk>
	`籠`: [u8(0xE2), 0xC4] // U+7C60 <cjk>
	`簀`: [u8(0xE2), 0xC5] // U+7C00 <cjk>
	`簇`: [u8(0xE2), 0xC6] // U+7C07 <cjk>
	`簓`: [u8(0xE2), 0xC7] // U+7C13 <cjk>
	`篳`: [u8(0xE2), 0xC8] // U+7BF3 <cjk>
	`篷`: [u8(0xE2), 0xC9] // U+7BF7 <cjk>
	`簗`: [u8(0xE2), 0xCA] // U+7C17 <cjk>
	`簍`: [u8(0xE2), 0xCB] // U+7C0D <cjk>
	`篶`: [u8(0xE2), 0xCC] // U+7BF6 <cjk>
	`簣`: [u8(0xE2), 0xCD] // U+7C23 <cjk>
	`簧`: [u8(0xE2), 0xCE] // U+7C27 <cjk>
	`簪`: [u8(0xE2), 0xCF] // U+7C2A <cjk>
	`簟`: [u8(0xE2), 0xD0] // U+7C1F <cjk>
	`簷`: [u8(0xE2), 0xD1] // U+7C37 <cjk>
	`簫`: [u8(0xE2), 0xD2] // U+7C2B <cjk>
	`簽`: [u8(0xE2), 0xD3] // U+7C3D <cjk>
	`籌`: [u8(0xE2), 0xD4] // U+7C4C <cjk>
	`籃`: [u8(0xE2), 0xD5] // U+7C43 <cjk>
	`籔`: [u8(0xE2), 0xD6] // U+7C54 <cjk>
	`籏`: [u8(0xE2), 0xD7] // U+7C4F <cjk>
	`籀`: [u8(0xE2), 0xD8] // U+7C40 <cjk>
	`籐`: [u8(0xE2), 0xD9] // U+7C50 <cjk>
	`籘`: [u8(0xE2), 0xDA] // U+7C58 <cjk>
	`籟`: [u8(0xE2), 0xDB] // U+7C5F <cjk>
	`籤`: [u8(0xE2), 0xDC] // U+7C64 <cjk>
	`籖`: [u8(0xE2), 0xDD] // U+7C56 <cjk>
	`籥`: [u8(0xE2), 0xDE] // U+7C65 <cjk>
	`籬`: [u8(0xE2), 0xDF] // U+7C6C <cjk>
	`籵`: [u8(0xE2), 0xE0] // U+7C75 <cjk>
	`粃`: [u8(0xE2), 0xE1] // U+7C83 <cjk>
	`粐`: [u8(0xE2), 0xE2] // U+7C90 <cjk>
	`粤`: [u8(0xE2), 0xE3] // U+7CA4 <cjk>
	`粭`: [u8(0xE2), 0xE4] // U+7CAD <cjk>
	`粢`: [u8(0xE2), 0xE5] // U+7CA2 <cjk>
	`粫`: [u8(0xE2), 0xE6] // U+7CAB <cjk>
	`粡`: [u8(0xE2), 0xE7] // U+7CA1 <cjk>
	`粨`: [u8(0xE2), 0xE8] // U+7CA8 <cjk>
	`粳`: [u8(0xE2), 0xE9] // U+7CB3 <cjk>
	`粲`: [u8(0xE2), 0xEA] // U+7CB2 <cjk>
	`粱`: [u8(0xE2), 0xEB] // U+7CB1 <cjk>
	`粮`: [u8(0xE2), 0xEC] // U+7CAE <cjk>
	`粹`: [u8(0xE2), 0xED] // U+7CB9 <cjk>
	`粽`: [u8(0xE2), 0xEE] // U+7CBD <cjk>
	`糀`: [u8(0xE2), 0xEF] // U+7CC0 <cjk>
	`糅`: [u8(0xE2), 0xF0] // U+7CC5 <cjk>
	`糂`: [u8(0xE2), 0xF1] // U+7CC2 <cjk>
	`糘`: [u8(0xE2), 0xF2] // U+7CD8 <cjk>
	`糒`: [u8(0xE2), 0xF3] // U+7CD2 <cjk>
	`糜`: [u8(0xE2), 0xF4] // U+7CDC <cjk>
	`糢`: [u8(0xE2), 0xF5] // U+7CE2 <cjk>
	`鬻`: [u8(0xE2), 0xF6] // U+9B3B <cjk>
	`糯`: [u8(0xE2), 0xF7] // U+7CEF <cjk>
	`糲`: [u8(0xE2), 0xF8] // U+7CF2 <cjk>
	`糴`: [u8(0xE2), 0xF9] // U+7CF4 <cjk>
	`糶`: [u8(0xE2), 0xFA] // U+7CF6 <cjk>
	`糺`: [u8(0xE2), 0xFB] // U+7CFA <cjk>
	`紆`: [u8(0xE2), 0xFC] // U+7D06 <cjk>
	`紂`: [u8(0xE3), 0x40] // U+7D02 <cjk>
	`紜`: [u8(0xE3), 0x41] // U+7D1C <cjk>
	`紕`: [u8(0xE3), 0x42] // U+7D15 <cjk>
	`紊`: [u8(0xE3), 0x43] // U+7D0A <cjk>
	`絅`: [u8(0xE3), 0x44] // U+7D45 <cjk>
	`絋`: [u8(0xE3), 0x45] // U+7D4B <cjk>
	`紮`: [u8(0xE3), 0x46] // U+7D2E <cjk>
	`紲`: [u8(0xE3), 0x47] // U+7D32 <cjk>
	`紿`: [u8(0xE3), 0x48] // U+7D3F <cjk>
	`紵`: [u8(0xE3), 0x49] // U+7D35 <cjk>
	`絆`: [u8(0xE3), 0x4A] // U+7D46 <cjk>
	`絳`: [u8(0xE3), 0x4B] // U+7D73 <cjk>
	`絖`: [u8(0xE3), 0x4C] // U+7D56 <cjk>
	`絎`: [u8(0xE3), 0x4D] // U+7D4E <cjk>
	`絲`: [u8(0xE3), 0x4E] // U+7D72 <cjk>
	`絨`: [u8(0xE3), 0x4F] // U+7D68 <cjk>
	`絮`: [u8(0xE3), 0x50] // U+7D6E <cjk>
	`絏`: [u8(0xE3), 0x51] // U+7D4F <cjk>
	`絣`: [u8(0xE3), 0x52] // U+7D63 <cjk>
	`經`: [u8(0xE3), 0x53] // U+7D93 <cjk>
	`綉`: [u8(0xE3), 0x54] // U+7D89 <cjk>
	`絛`: [u8(0xE3), 0x55] // U+7D5B <cjk>
	`綏`: [u8(0xE3), 0x56] // U+7D8F <cjk>
	`絽`: [u8(0xE3), 0x57] // U+7D7D <cjk>
	`綛`: [u8(0xE3), 0x58] // U+7D9B <cjk>
	`綺`: [u8(0xE3), 0x59] // U+7DBA <cjk>
	`綮`: [u8(0xE3), 0x5A] // U+7DAE <cjk>
	`綣`: [u8(0xE3), 0x5B] // U+7DA3 <cjk>
	`綵`: [u8(0xE3), 0x5C] // U+7DB5 <cjk>
	`緇`: [u8(0xE3), 0x5D] // U+7DC7 <cjk>
	`綽`: [u8(0xE3), 0x5E] // U+7DBD <cjk>
	`綫`: [u8(0xE3), 0x5F] // U+7DAB <cjk>
	`總`: [u8(0xE3), 0x60] // U+7E3D <cjk>
	`綢`: [u8(0xE3), 0x61] // U+7DA2 <cjk>
	`綯`: [u8(0xE3), 0x62] // U+7DAF <cjk>
	`緜`: [u8(0xE3), 0x63] // U+7DDC <cjk>
	`綸`: [u8(0xE3), 0x64] // U+7DB8 <cjk>
	`綟`: [u8(0xE3), 0x65] // U+7D9F <cjk>
	`綰`: [u8(0xE3), 0x66] // U+7DB0 <cjk>
	`緘`: [u8(0xE3), 0x67] // U+7DD8 <cjk>
	`緝`: [u8(0xE3), 0x68] // U+7DDD <cjk>
	`緤`: [u8(0xE3), 0x69] // U+7DE4 <cjk>
	`緞`: [u8(0xE3), 0x6A] // U+7DDE <cjk>
	`緻`: [u8(0xE3), 0x6B] // U+7DFB <cjk>
	`緲`: [u8(0xE3), 0x6C] // U+7DF2 <cjk>
	`緡`: [u8(0xE3), 0x6D] // U+7DE1 <cjk>
	`縅`: [u8(0xE3), 0x6E] // U+7E05 <cjk>
	`縊`: [u8(0xE3), 0x6F] // U+7E0A <cjk>
	`縣`: [u8(0xE3), 0x70] // U+7E23 <cjk>
	`縡`: [u8(0xE3), 0x71] // U+7E21 <cjk>
	`縒`: [u8(0xE3), 0x72] // U+7E12 <cjk>
	`縱`: [u8(0xE3), 0x73] // U+7E31 <cjk>
	`縟`: [u8(0xE3), 0x74] // U+7E1F <cjk>
	`縉`: [u8(0xE3), 0x75] // U+7E09 <cjk>
	`縋`: [u8(0xE3), 0x76] // U+7E0B <cjk>
	`縢`: [u8(0xE3), 0x77] // U+7E22 <cjk>
	`繆`: [u8(0xE3), 0x78] // U+7E46 <cjk>
	`繦`: [u8(0xE3), 0x79] // U+7E66 <cjk>
	`縻`: [u8(0xE3), 0x7A] // U+7E3B <cjk>
	`縵`: [u8(0xE3), 0x7B] // U+7E35 <cjk>
	`縹`: [u8(0xE3), 0x7C] // U+7E39 <cjk>
	`繃`: [u8(0xE3), 0x7D] // U+7E43 <cjk>
	`縷`: [u8(0xE3), 0x7E] // U+7E37 <cjk>
	`縲`: [u8(0xE3), 0x80] // U+7E32 <cjk>
	`縺`: [u8(0xE3), 0x81] // U+7E3A <cjk>
	`繧`: [u8(0xE3), 0x82] // U+7E67 <cjk>
	`繝`: [u8(0xE3), 0x83] // U+7E5D <cjk>
	`繖`: [u8(0xE3), 0x84] // U+7E56 <cjk>
	`繞`: [u8(0xE3), 0x85] // U+7E5E <cjk>
	`繙`: [u8(0xE3), 0x86] // U+7E59 <cjk>
	`繚`: [u8(0xE3), 0x87] // U+7E5A <cjk>
	`繹`: [u8(0xE3), 0x88] // U+7E79 <cjk>
	`繪`: [u8(0xE3), 0x89] // U+7E6A <cjk>
	`繩`: [u8(0xE3), 0x8A] // U+7E69 <cjk>
	`繼`: [u8(0xE3), 0x8B] // U+7E7C <cjk>
	`繻`: [u8(0xE3), 0x8C] // U+7E7B <cjk>
	`纃`: [u8(0xE3), 0x8D] // U+7E83 <cjk>
	`緕`: [u8(0xE3), 0x8E] // U+7DD5 <cjk>
	`繽`: [u8(0xE3), 0x8F] // U+7E7D <cjk>
	`辮`: [u8(0xE3), 0x90] // U+8FAE <cjk>
	`繿`: [u8(0xE3), 0x91] // U+7E7F <cjk>
	`纈`: [u8(0xE3), 0x92] // U+7E88 <cjk>
	`纉`: [u8(0xE3), 0x93] // U+7E89 <cjk>
	`續`: [u8(0xE3), 0x94] // U+7E8C <cjk>
	`纒`: [u8(0xE3), 0x95] // U+7E92 <cjk>
	`纐`: [u8(0xE3), 0x96] // U+7E90 <cjk>
	`纓`: [u8(0xE3), 0x97] // U+7E93 <cjk>
	`纔`: [u8(0xE3), 0x98] // U+7E94 <cjk>
	`纖`: [u8(0xE3), 0x99] // U+7E96 <cjk>
	`纎`: [u8(0xE3), 0x9A] // U+7E8E <cjk>
	`纛`: [u8(0xE3), 0x9B] // U+7E9B <cjk>
	`纜`: [u8(0xE3), 0x9C] // U+7E9C <cjk>
	`缸`: [u8(0xE3), 0x9D] // U+7F38 <cjk>
	`缺`: [u8(0xE3), 0x9E] // U+7F3A <cjk>
	`罅`: [u8(0xE3), 0x9F] // U+7F45 <cjk>
	`罌`: [u8(0xE3), 0xA0] // U+7F4C <cjk>
	`罍`: [u8(0xE3), 0xA1] // U+7F4D <cjk>
	`罎`: [u8(0xE3), 0xA2] // U+7F4E <cjk>
	`罐`: [u8(0xE3), 0xA3] // U+7F50 <cjk>
	`网`: [u8(0xE3), 0xA4] // U+7F51 <cjk>
	`罕`: [u8(0xE3), 0xA5] // U+7F55 <cjk>
	`罔`: [u8(0xE3), 0xA6] // U+7F54 <cjk>
	`罘`: [u8(0xE3), 0xA7] // U+7F58 <cjk>
	`罟`: [u8(0xE3), 0xA8] // U+7F5F <cjk>
	`罠`: [u8(0xE3), 0xA9] // U+7F60 <cjk>
	`罨`: [u8(0xE3), 0xAA] // U+7F68 <cjk>
	`罩`: [u8(0xE3), 0xAB] // U+7F69 <cjk>
	`罧`: [u8(0xE3), 0xAC] // U+7F67 <cjk>
	`罸`: [u8(0xE3), 0xAD] // U+7F78 <cjk>
	`羂`: [u8(0xE3), 0xAE] // U+7F82 <cjk>
	`羆`: [u8(0xE3), 0xAF] // U+7F86 <cjk>
	`羃`: [u8(0xE3), 0xB0] // U+7F83 <cjk>
	`羈`: [u8(0xE3), 0xB1] // U+7F88 <cjk>
	`羇`: [u8(0xE3), 0xB2] // U+7F87 <cjk>
	`羌`: [u8(0xE3), 0xB3] // U+7F8C <cjk>
	`羔`: [u8(0xE3), 0xB4] // U+7F94 <cjk>
	`羞`: [u8(0xE3), 0xB5] // U+7F9E <cjk>
	`羝`: [u8(0xE3), 0xB6] // U+7F9D <cjk>
	`羚`: [u8(0xE3), 0xB7] // U+7F9A <cjk>
	`羣`: [u8(0xE3), 0xB8] // U+7FA3 <cjk>
	`羯`: [u8(0xE3), 0xB9] // U+7FAF <cjk>
	`羲`: [u8(0xE3), 0xBA] // U+7FB2 <cjk>
	`羹`: [u8(0xE3), 0xBB] // U+7FB9 <cjk>
	`羮`: [u8(0xE3), 0xBC] // U+7FAE <cjk>
	`羶`: [u8(0xE3), 0xBD] // U+7FB6 <cjk>
	`羸`: [u8(0xE3), 0xBE] // U+7FB8 <cjk>
	`譱`: [u8(0xE3), 0xBF] // U+8B71 <cjk>
	`翅`: [u8(0xE3), 0xC0] // U+7FC5 <cjk>
	`翆`: [u8(0xE3), 0xC1] // U+7FC6 <cjk>
	`翊`: [u8(0xE3), 0xC2] // U+7FCA <cjk>
	`翕`: [u8(0xE3), 0xC3] // U+7FD5 <cjk>
	`翔`: [u8(0xE3), 0xC4] // U+7FD4 <cjk>
	`翡`: [u8(0xE3), 0xC5] // U+7FE1 <cjk>
	`翦`: [u8(0xE3), 0xC6] // U+7FE6 <cjk>
	`翩`: [u8(0xE3), 0xC7] // U+7FE9 <cjk>
	`翳`: [u8(0xE3), 0xC8] // U+7FF3 <cjk>
	`翹`: [u8(0xE3), 0xC9] // U+7FF9 <cjk>
	`飜`: [u8(0xE3), 0xCA] // U+98DC <cjk>
	`耆`: [u8(0xE3), 0xCB] // U+8006 <cjk>
	`耄`: [u8(0xE3), 0xCC] // U+8004 <cjk>
	`耋`: [u8(0xE3), 0xCD] // U+800B <cjk>
	`耒`: [u8(0xE3), 0xCE] // U+8012 <cjk>
	`耘`: [u8(0xE3), 0xCF] // U+8018 <cjk>
	`耙`: [u8(0xE3), 0xD0] // U+8019 <cjk>
	`耜`: [u8(0xE3), 0xD1] // U+801C <cjk>
	`耡`: [u8(0xE3), 0xD2] // U+8021 <cjk>
	`耨`: [u8(0xE3), 0xD3] // U+8028 <cjk>
	`耿`: [u8(0xE3), 0xD4] // U+803F <cjk>
	`耻`: [u8(0xE3), 0xD5] // U+803B <cjk>
	`聊`: [u8(0xE3), 0xD6] // U+804A <cjk>
	`聆`: [u8(0xE3), 0xD7] // U+8046 <cjk>
	`聒`: [u8(0xE3), 0xD8] // U+8052 <cjk>
	`聘`: [u8(0xE3), 0xD9] // U+8058 <cjk>
	`聚`: [u8(0xE3), 0xDA] // U+805A <cjk>
	`聟`: [u8(0xE3), 0xDB] // U+805F <cjk>
	`聢`: [u8(0xE3), 0xDC] // U+8062 <cjk>
	`聨`: [u8(0xE3), 0xDD] // U+8068 <cjk>
	`聳`: [u8(0xE3), 0xDE] // U+8073 <cjk>
	`聲`: [u8(0xE3), 0xDF] // U+8072 <cjk>
	`聰`: [u8(0xE3), 0xE0] // U+8070 <cjk>
	`聶`: [u8(0xE3), 0xE1] // U+8076 <cjk>
	`聹`: [u8(0xE3), 0xE2] // U+8079 <cjk>
	`聽`: [u8(0xE3), 0xE3] // U+807D <cjk>
	`聿`: [u8(0xE3), 0xE4] // U+807F <cjk>
	`肄`: [u8(0xE3), 0xE5] // U+8084 <cjk>
	`肆`: [u8(0xE3), 0xE6] // U+8086 <cjk>
	`肅`: [u8(0xE3), 0xE7] // U+8085 <cjk>
	`肛`: [u8(0xE3), 0xE8] // U+809B <cjk>
	`肓`: [u8(0xE3), 0xE9] // U+8093 <cjk>
	`肚`: [u8(0xE3), 0xEA] // U+809A <cjk>
	`肭`: [u8(0xE3), 0xEB] // U+80AD <cjk>
	`冐`: [u8(0xE3), 0xEC] // U+5190 <cjk>
	`肬`: [u8(0xE3), 0xED] // U+80AC <cjk>
	`胛`: [u8(0xE3), 0xEE] // U+80DB <cjk>
	`胥`: [u8(0xE3), 0xEF] // U+80E5 <cjk>
	`胙`: [u8(0xE3), 0xF0] // U+80D9 <cjk>
	`胝`: [u8(0xE3), 0xF1] // U+80DD <cjk>
	`胄`: [u8(0xE3), 0xF2] // U+80C4 <cjk>
	`胚`: [u8(0xE3), 0xF3] // U+80DA <cjk>
	`胖`: [u8(0xE3), 0xF4] // U+80D6 <cjk>
	`脉`: [u8(0xE3), 0xF5] // U+8109 <cjk>
	`胯`: [u8(0xE3), 0xF6] // U+80EF <cjk>
	`胱`: [u8(0xE3), 0xF7] // U+80F1 <cjk>
	`脛`: [u8(0xE3), 0xF8] // U+811B <cjk>
	`脩`: [u8(0xE3), 0xF9] // U+8129 <cjk>
	`脣`: [u8(0xE3), 0xFA] // U+8123 <cjk>
	`脯`: [u8(0xE3), 0xFB] // U+812F <cjk>
	`腋`: [u8(0xE3), 0xFC] // U+814B <cjk>
	`隋`: [u8(0xE4), 0x40] // U+968B <cjk>
	`腆`: [u8(0xE4), 0x41] // U+8146 <cjk>
	`脾`: [u8(0xE4), 0x42] // U+813E <cjk>
	`腓`: [u8(0xE4), 0x43] // U+8153 <cjk>
	`腑`: [u8(0xE4), 0x44] // U+8151 <cjk>
	`胼`: [u8(0xE4), 0x45] // U+80FC <cjk>
	`腱`: [u8(0xE4), 0x46] // U+8171 <cjk>
	`腮`: [u8(0xE4), 0x47] // U+816E <cjk>
	`腥`: [u8(0xE4), 0x48] // U+8165 <cjk>
	`腦`: [u8(0xE4), 0x49] // U+8166 <cjk>
	`腴`: [u8(0xE4), 0x4A] // U+8174 <cjk>
	`膃`: [u8(0xE4), 0x4B] // U+8183 <cjk>
	`膈`: [u8(0xE4), 0x4C] // U+8188 <cjk>
	`膊`: [u8(0xE4), 0x4D] // U+818A <cjk>
	`膀`: [u8(0xE4), 0x4E] // U+8180 <cjk>
	`膂`: [u8(0xE4), 0x4F] // U+8182 <cjk>
	`膠`: [u8(0xE4), 0x50] // U+81A0 <cjk>
	`膕`: [u8(0xE4), 0x51] // U+8195 <cjk>
	`膤`: [u8(0xE4), 0x52] // U+81A4 <cjk>
	`膣`: [u8(0xE4), 0x53] // U+81A3 <cjk>
	`腟`: [u8(0xE4), 0x54] // U+815F <cjk>
	`膓`: [u8(0xE4), 0x55] // U+8193 <cjk>
	`膩`: [u8(0xE4), 0x56] // U+81A9 <cjk>
	`膰`: [u8(0xE4), 0x57] // U+81B0 <cjk>
	`膵`: [u8(0xE4), 0x58] // U+81B5 <cjk>
	`膾`: [u8(0xE4), 0x59] // U+81BE <cjk>
	`膸`: [u8(0xE4), 0x5A] // U+81B8 <cjk>
	`膽`: [u8(0xE4), 0x5B] // U+81BD <cjk>
	`臀`: [u8(0xE4), 0x5C] // U+81C0 <cjk>
	`臂`: [u8(0xE4), 0x5D] // U+81C2 <cjk>
	`膺`: [u8(0xE4), 0x5E] // U+81BA <cjk>
	`臉`: [u8(0xE4), 0x5F] // U+81C9 <cjk>
	`臍`: [u8(0xE4), 0x60] // U+81CD <cjk>
	`臑`: [u8(0xE4), 0x61] // U+81D1 <cjk>
	`臙`: [u8(0xE4), 0x62] // U+81D9 <cjk>
	`臘`: [u8(0xE4), 0x63] // U+81D8 <cjk>
	`臈`: [u8(0xE4), 0x64] // U+81C8 <cjk>
	`臚`: [u8(0xE4), 0x65] // U+81DA <cjk>
	`臟`: [u8(0xE4), 0x66] // U+81DF <cjk>
	`臠`: [u8(0xE4), 0x67] // U+81E0 <cjk>
	`臧`: [u8(0xE4), 0x68] // U+81E7 <cjk>
	`臺`: [u8(0xE4), 0x69] // U+81FA <cjk>
	`臻`: [u8(0xE4), 0x6A] // U+81FB <cjk>
	`臾`: [u8(0xE4), 0x6B] // U+81FE <cjk>
	`舁`: [u8(0xE4), 0x6C] // U+8201 <cjk>
	`舂`: [u8(0xE4), 0x6D] // U+8202 <cjk>
	`舅`: [u8(0xE4), 0x6E] // U+8205 <cjk>
	`與`: [u8(0xE4), 0x6F] // U+8207 <cjk>
	`舊`: [u8(0xE4), 0x70] // U+820A <cjk>
	`舍`: [u8(0xE4), 0x71] // U+820D <cjk>
	`舐`: [u8(0xE4), 0x72] // U+8210 <cjk>
	`舖`: [u8(0xE4), 0x73] // U+8216 <cjk>
	`舩`: [u8(0xE4), 0x74] // U+8229 <cjk>
	`舫`: [u8(0xE4), 0x75] // U+822B <cjk>
	`舸`: [u8(0xE4), 0x76] // U+8238 <cjk>
	`舳`: [u8(0xE4), 0x77] // U+8233 <cjk>
	`艀`: [u8(0xE4), 0x78] // U+8240 <cjk>
	`艙`: [u8(0xE4), 0x79] // U+8259 <cjk>
	`艘`: [u8(0xE4), 0x7A] // U+8258 <cjk>
	`艝`: [u8(0xE4), 0x7B] // U+825D <cjk>
	`艚`: [u8(0xE4), 0x7C] // U+825A <cjk>
	`艟`: [u8(0xE4), 0x7D] // U+825F <cjk>
	`艤`: [u8(0xE4), 0x7E] // U+8264 <cjk>
	`艢`: [u8(0xE4), 0x80] // U+8262 <cjk>
	`艨`: [u8(0xE4), 0x81] // U+8268 <cjk>
	`艪`: [u8(0xE4), 0x82] // U+826A <cjk>
	`艫`: [u8(0xE4), 0x83] // U+826B <cjk>
	`舮`: [u8(0xE4), 0x84] // U+822E <cjk>
	`艱`: [u8(0xE4), 0x85] // U+8271 <cjk>
	`艷`: [u8(0xE4), 0x86] // U+8277 <cjk>
	`艸`: [u8(0xE4), 0x87] // U+8278 <cjk>
	`艾`: [u8(0xE4), 0x88] // U+827E <cjk>
	`芍`: [u8(0xE4), 0x89] // U+828D <cjk>
	`芒`: [u8(0xE4), 0x8A] // U+8292 <cjk>
	`芫`: [u8(0xE4), 0x8B] // U+82AB <cjk>
	`芟`: [u8(0xE4), 0x8C] // U+829F <cjk>
	`芻`: [u8(0xE4), 0x8D] // U+82BB <cjk>
	`芬`: [u8(0xE4), 0x8E] // U+82AC <cjk>
	`苡`: [u8(0xE4), 0x8F] // U+82E1 <cjk>
	`苣`: [u8(0xE4), 0x90] // U+82E3 <cjk>
	`苟`: [u8(0xE4), 0x91] // U+82DF <cjk>
	`苒`: [u8(0xE4), 0x92] // U+82D2 <cjk>
	`苴`: [u8(0xE4), 0x93] // U+82F4 <cjk>
	`苳`: [u8(0xE4), 0x94] // U+82F3 <cjk>
	`苺`: [u8(0xE4), 0x95] // U+82FA <cjk>
	`莓`: [u8(0xE4), 0x96] // U+8393 <cjk>
	`范`: [u8(0xE4), 0x97] // U+8303 <cjk>
	`苻`: [u8(0xE4), 0x98] // U+82FB <cjk>
	`苹`: [u8(0xE4), 0x99] // U+82F9 <cjk>
	`苞`: [u8(0xE4), 0x9A] // U+82DE <cjk>
	`茆`: [u8(0xE4), 0x9B] // U+8306 <cjk>
	`苜`: [u8(0xE4), 0x9C] // U+82DC <cjk>
	`茉`: [u8(0xE4), 0x9D] // U+8309 <cjk>
	`苙`: [u8(0xE4), 0x9E] // U+82D9 <cjk>
	`茵`: [u8(0xE4), 0x9F] // U+8335 <cjk>
	`茴`: [u8(0xE4), 0xA0] // U+8334 <cjk>
	`茖`: [u8(0xE4), 0xA1] // U+8316 <cjk>
	`茲`: [u8(0xE4), 0xA2] // U+8332 <cjk>
	`茱`: [u8(0xE4), 0xA3] // U+8331 <cjk>
	`荀`: [u8(0xE4), 0xA4] // U+8340 <cjk>
	`茹`: [u8(0xE4), 0xA5] // U+8339 <cjk>
	`荐`: [u8(0xE4), 0xA6] // U+8350 <cjk>
	`荅`: [u8(0xE4), 0xA7] // U+8345 <cjk>
	`茯`: [u8(0xE4), 0xA8] // U+832F <cjk>
	`茫`: [u8(0xE4), 0xA9] // U+832B <cjk>
	`茗`: [u8(0xE4), 0xAA] // U+8317 <cjk>
	`茘`: [u8(0xE4), 0xAB] // U+8318 <cjk>
	`莅`: [u8(0xE4), 0xAC] // U+8385 <cjk>
	`莚`: [u8(0xE4), 0xAD] // U+839A <cjk>
	`莪`: [u8(0xE4), 0xAE] // U+83AA <cjk>
	`莟`: [u8(0xE4), 0xAF] // U+839F <cjk>
	`莢`: [u8(0xE4), 0xB0] // U+83A2 <cjk>
	`莖`: [u8(0xE4), 0xB1] // U+8396 <cjk>
	`茣`: [u8(0xE4), 0xB2] // U+8323 <cjk>
	`莎`: [u8(0xE4), 0xB3] // U+838E <cjk>
	`莇`: [u8(0xE4), 0xB4] // U+8387 <cjk>
	`莊`: [u8(0xE4), 0xB5] // U+838A <cjk>
	`荼`: [u8(0xE4), 0xB6] // U+837C <cjk>
	`莵`: [u8(0xE4), 0xB7] // U+83B5 <cjk>
	`荳`: [u8(0xE4), 0xB8] // U+8373 <cjk>
	`荵`: [u8(0xE4), 0xB9] // U+8375 <cjk>
	`莠`: [u8(0xE4), 0xBA] // U+83A0 <cjk>
	`莉`: [u8(0xE4), 0xBB] // U+8389 <cjk>
	`莨`: [u8(0xE4), 0xBC] // U+83A8 <cjk>
	`菴`: [u8(0xE4), 0xBD] // U+83F4 <cjk>
	`萓`: [u8(0xE4), 0xBE] // U+8413 <cjk>
	`菫`: [u8(0xE4), 0xBF] // U+83EB <cjk>
	`菎`: [u8(0xE4), 0xC0] // U+83CE <cjk>
	`菽`: [u8(0xE4), 0xC1] // U+83FD <cjk>
	`萃`: [u8(0xE4), 0xC2] // U+8403 <cjk>
	`菘`: [u8(0xE4), 0xC3] // U+83D8 <cjk>
	`萋`: [u8(0xE4), 0xC4] // U+840B <cjk>
	`菁`: [u8(0xE4), 0xC5] // U+83C1 <cjk>
	`菷`: [u8(0xE4), 0xC6] // U+83F7 <cjk>
	`萇`: [u8(0xE4), 0xC7] // U+8407 <cjk>
	`菠`: [u8(0xE4), 0xC8] // U+83E0 <cjk>
	`菲`: [u8(0xE4), 0xC9] // U+83F2 <cjk>
	`萍`: [u8(0xE4), 0xCA] // U+840D <cjk>
	`萢`: [u8(0xE4), 0xCB] // U+8422 <cjk>
	`萠`: [u8(0xE4), 0xCC] // U+8420 <cjk>
	`莽`: [u8(0xE4), 0xCD] // U+83BD <cjk>
	`萸`: [u8(0xE4), 0xCE] // U+8438 <cjk>
	`蔆`: [u8(0xE4), 0xCF] // U+8506 <cjk>
	`菻`: [u8(0xE4), 0xD0] // U+83FB <cjk>
	`葭`: [u8(0xE4), 0xD1] // U+846D <cjk>
	`萪`: [u8(0xE4), 0xD2] // U+842A <cjk>
	`萼`: [u8(0xE4), 0xD3] // U+843C <cjk>
	`蕚`: [u8(0xE4), 0xD4] // U+855A <cjk>
	`蒄`: [u8(0xE4), 0xD5] // U+8484 <cjk>
	`葷`: [u8(0xE4), 0xD6] // U+8477 <cjk>
	`葫`: [u8(0xE4), 0xD7] // U+846B <cjk>
	`蒭`: [u8(0xE4), 0xD8] // U+84AD <cjk>
	`葮`: [u8(0xE4), 0xD9] // U+846E <cjk>
	`蒂`: [u8(0xE4), 0xDA] // U+8482 <cjk>
	`葩`: [u8(0xE4), 0xDB] // U+8469 <cjk>
	`葆`: [u8(0xE4), 0xDC] // U+8446 <cjk>
	`萬`: [u8(0xE4), 0xDD] // U+842C <cjk>
	`葯`: [u8(0xE4), 0xDE] // U+846F <cjk>
	`葹`: [u8(0xE4), 0xDF] // U+8479 <cjk>
	`萵`: [u8(0xE4), 0xE0] // U+8435 <cjk>
	`蓊`: [u8(0xE4), 0xE1] // U+84CA <cjk>
	`葢`: [u8(0xE4), 0xE2] // U+8462 <cjk>
	`蒹`: [u8(0xE4), 0xE3] // U+84B9 <cjk>
	`蒿`: [u8(0xE4), 0xE4] // U+84BF <cjk>
	`蒟`: [u8(0xE4), 0xE5] // U+849F <cjk>
	`蓙`: [u8(0xE4), 0xE6] // U+84D9 <cjk>
	`蓍`: [u8(0xE4), 0xE7] // U+84CD <cjk>
	`蒻`: [u8(0xE4), 0xE8] // U+84BB <cjk>
	`蓚`: [u8(0xE4), 0xE9] // U+84DA <cjk>
	`蓐`: [u8(0xE4), 0xEA] // U+84D0 <cjk>
	`蓁`: [u8(0xE4), 0xEB] // U+84C1 <cjk>
	`蓆`: [u8(0xE4), 0xEC] // U+84C6 <cjk>
	`蓖`: [u8(0xE4), 0xED] // U+84D6 <cjk>
	`蒡`: [u8(0xE4), 0xEE] // U+84A1 <cjk>
	`蔡`: [u8(0xE4), 0xEF] // U+8521 <cjk>
	`蓿`: [u8(0xE4), 0xF0] // U+84FF <cjk>
	`蓴`: [u8(0xE4), 0xF1] // U+84F4 <cjk>
	`蔗`: [u8(0xE4), 0xF2] // U+8517 <cjk>
	`蔘`: [u8(0xE4), 0xF3] // U+8518 <cjk>
	`蔬`: [u8(0xE4), 0xF4] // U+852C <cjk>
	`蔟`: [u8(0xE4), 0xF5] // U+851F <cjk>
	`蔕`: [u8(0xE4), 0xF6] // U+8515 <cjk>
	`蔔`: [u8(0xE4), 0xF7] // U+8514 <cjk>
	`蓼`: [u8(0xE4), 0xF8] // U+84FC <cjk>
	`蕀`: [u8(0xE4), 0xF9] // U+8540 <cjk>
	`蕣`: [u8(0xE4), 0xFA] // U+8563 <cjk>
	`蕘`: [u8(0xE4), 0xFB] // U+8558 <cjk>
	`蕈`: [u8(0xE4), 0xFC] // U+8548 <cjk>
	`蕁`: [u8(0xE5), 0x40] // U+8541 <cjk>
	`蘂`: [u8(0xE5), 0x41] // U+8602 <cjk>
	`蕋`: [u8(0xE5), 0x42] // U+854B <cjk>
	`蕕`: [u8(0xE5), 0x43] // U+8555 <cjk>
	`薀`: [u8(0xE5), 0x44] // U+8580 <cjk>
	`薤`: [u8(0xE5), 0x45] // U+85A4 <cjk>
	`薈`: [u8(0xE5), 0x46] // U+8588 <cjk>
	`薑`: [u8(0xE5), 0x47] // U+8591 <cjk>
	`薊`: [u8(0xE5), 0x48] // U+858A <cjk>
	`薨`: [u8(0xE5), 0x49] // U+85A8 <cjk>
	`蕭`: [u8(0xE5), 0x4A] // U+856D <cjk>
	`薔`: [u8(0xE5), 0x4B] // U+8594 <cjk>
	`薛`: [u8(0xE5), 0x4C] // U+859B <cjk>
	`藪`: [u8(0xE5), 0x4D] // U+85EA <cjk>
	`薇`: [u8(0xE5), 0x4E] // U+8587 <cjk>
	`薜`: [u8(0xE5), 0x4F] // U+859C <cjk>
	`蕷`: [u8(0xE5), 0x50] // U+8577 <cjk>
	`蕾`: [u8(0xE5), 0x51] // U+857E <cjk>
	`薐`: [u8(0xE5), 0x52] // U+8590 <cjk>
	`藉`: [u8(0xE5), 0x53] // U+85C9 <cjk>
	`薺`: [u8(0xE5), 0x54] // U+85BA <cjk>
	`藏`: [u8(0xE5), 0x55] // U+85CF <cjk>
	`薹`: [u8(0xE5), 0x56] // U+85B9 <cjk>
	`藐`: [u8(0xE5), 0x57] // U+85D0 <cjk>
	`藕`: [u8(0xE5), 0x58] // U+85D5 <cjk>
	`藝`: [u8(0xE5), 0x59] // U+85DD <cjk>
	`藥`: [u8(0xE5), 0x5A] // U+85E5 <cjk>
	`藜`: [u8(0xE5), 0x5B] // U+85DC <cjk>
	`藹`: [u8(0xE5), 0x5C] // U+85F9 <cjk>
	`蘊`: [u8(0xE5), 0x5D] // U+860A <cjk>
	`蘓`: [u8(0xE5), 0x5E] // U+8613 <cjk>
	`蘋`: [u8(0xE5), 0x5F] // U+860B <cjk>
	`藾`: [u8(0xE5), 0x60] // U+85FE <cjk>
	`藺`: [u8(0xE5), 0x61] // U+85FA <cjk>
	`蘆`: [u8(0xE5), 0x62] // U+8606 <cjk>
	`蘢`: [u8(0xE5), 0x63] // U+8622 <cjk>
	`蘚`: [u8(0xE5), 0x64] // U+861A <cjk>
	`蘰`: [u8(0xE5), 0x65] // U+8630 <cjk>
	`蘿`: [u8(0xE5), 0x66] // U+863F <cjk>
	`虍`: [u8(0xE5), 0x67] // U+864D <cjk>
	`乕`: [u8(0xE5), 0x68] // U+4E55 <cjk>
	`虔`: [u8(0xE5), 0x69] // U+8654 <cjk>
	`號`: [u8(0xE5), 0x6A] // U+865F <cjk>
	`虧`: [u8(0xE5), 0x6B] // U+8667 <cjk>
	`虱`: [u8(0xE5), 0x6C] // U+8671 <cjk>
	`蚓`: [u8(0xE5), 0x6D] // U+8693 <cjk>
	`蚣`: [u8(0xE5), 0x6E] // U+86A3 <cjk>
	`蚩`: [u8(0xE5), 0x6F] // U+86A9 <cjk>
	`蚪`: [u8(0xE5), 0x70] // U+86AA <cjk>
	`蚋`: [u8(0xE5), 0x71] // U+868B <cjk>
	`蚌`: [u8(0xE5), 0x72] // U+868C <cjk>
	`蚶`: [u8(0xE5), 0x73] // U+86B6 <cjk>
	`蚯`: [u8(0xE5), 0x74] // U+86AF <cjk>
	`蛄`: [u8(0xE5), 0x75] // U+86C4 <cjk>
	`蛆`: [u8(0xE5), 0x76] // U+86C6 <cjk>
	`蚰`: [u8(0xE5), 0x77] // U+86B0 <cjk>
	`蛉`: [u8(0xE5), 0x78] // U+86C9 <cjk>
	`蠣`: [u8(0xE5), 0x79] // U+8823 <cjk>
	`蚫`: [u8(0xE5), 0x7A] // U+86AB <cjk>
	`蛔`: [u8(0xE5), 0x7B] // U+86D4 <cjk>
	`蛞`: [u8(0xE5), 0x7C] // U+86DE <cjk>
	`蛩`: [u8(0xE5), 0x7D] // U+86E9 <cjk>
	`蛬`: [u8(0xE5), 0x7E] // U+86EC <cjk>
	`蛟`: [u8(0xE5), 0x80] // U+86DF <cjk>
	`蛛`: [u8(0xE5), 0x81] // U+86DB <cjk>
	`蛯`: [u8(0xE5), 0x82] // U+86EF <cjk>
	`蜒`: [u8(0xE5), 0x83] // U+8712 <cjk>
	`蜆`: [u8(0xE5), 0x84] // U+8706 <cjk>
	`蜈`: [u8(0xE5), 0x85] // U+8708 <cjk>
	`蜀`: [u8(0xE5), 0x86] // U+8700 <cjk>
	`蜃`: [u8(0xE5), 0x87] // U+8703 <cjk>
	`蛻`: [u8(0xE5), 0x88] // U+86FB <cjk>
	`蜑`: [u8(0xE5), 0x89] // U+8711 <cjk>
	`蜉`: [u8(0xE5), 0x8A] // U+8709 <cjk>
	`蜍`: [u8(0xE5), 0x8B] // U+870D <cjk>
	`蛹`: [u8(0xE5), 0x8C] // U+86F9 <cjk>
	`蜊`: [u8(0xE5), 0x8D] // U+870A <cjk>
	`蜴`: [u8(0xE5), 0x8E] // U+8734 <cjk>
	`蜿`: [u8(0xE5), 0x8F] // U+873F <cjk>
	`蜷`: [u8(0xE5), 0x90] // U+8737 <cjk>
	`蜻`: [u8(0xE5), 0x91] // U+873B <cjk>
	`蜥`: [u8(0xE5), 0x92] // U+8725 <cjk>
	`蜩`: [u8(0xE5), 0x93] // U+8729 <cjk>
	`蜚`: [u8(0xE5), 0x94] // U+871A <cjk>
	`蝠`: [u8(0xE5), 0x95] // U+8760 <cjk>
	`蝟`: [u8(0xE5), 0x96] // U+875F <cjk>
	`蝸`: [u8(0xE5), 0x97] // U+8778 <cjk>
	`蝌`: [u8(0xE5), 0x98] // U+874C <cjk>
	`蝎`: [u8(0xE5), 0x99] // U+874E <cjk>
	`蝴`: [u8(0xE5), 0x9A] // U+8774 <cjk>
	`蝗`: [u8(0xE5), 0x9B] // U+8757 <cjk>
	`蝨`: [u8(0xE5), 0x9C] // U+8768 <cjk>
	`蝮`: [u8(0xE5), 0x9D] // U+876E <cjk>
	`蝙`: [u8(0xE5), 0x9E] // U+8759 <cjk>
	`蝓`: [u8(0xE5), 0x9F] // U+8753 <cjk>
	`蝣`: [u8(0xE5), 0xA0] // U+8763 <cjk>
	`蝪`: [u8(0xE5), 0xA1] // U+876A <cjk>
	`蠅`: [u8(0xE5), 0xA2] // U+8805 <cjk>
	`螢`: [u8(0xE5), 0xA3] // U+87A2 <cjk>
	`螟`: [u8(0xE5), 0xA4] // U+879F <cjk>
	`螂`: [u8(0xE5), 0xA5] // U+8782 <cjk>
	`螯`: [u8(0xE5), 0xA6] // U+87AF <cjk>
	`蟋`: [u8(0xE5), 0xA7] // U+87CB <cjk>
	`螽`: [u8(0xE5), 0xA8] // U+87BD <cjk>
	`蟀`: [u8(0xE5), 0xA9] // U+87C0 <cjk>
	`蟐`: [u8(0xE5), 0xAA] // U+87D0 <cjk>
	`雖`: [u8(0xE5), 0xAB] // U+96D6 <cjk>
	`螫`: [u8(0xE5), 0xAC] // U+87AB <cjk>
	`蟄`: [u8(0xE5), 0xAD] // U+87C4 <cjk>
	`螳`: [u8(0xE5), 0xAE] // U+87B3 <cjk>
	`蟇`: [u8(0xE5), 0xAF] // U+87C7 <cjk>
	`蟆`: [u8(0xE5), 0xB0] // U+87C6 <cjk>
	`螻`: [u8(0xE5), 0xB1] // U+87BB <cjk>
	`蟯`: [u8(0xE5), 0xB2] // U+87EF <cjk>
	`蟲`: [u8(0xE5), 0xB3] // U+87F2 <cjk>
	`蟠`: [u8(0xE5), 0xB4] // U+87E0 <cjk>
	`蠏`: [u8(0xE5), 0xB5] // U+880F <cjk>
	`蠍`: [u8(0xE5), 0xB6] // U+880D <cjk>
	`蟾`: [u8(0xE5), 0xB7] // U+87FE <cjk>
	`蟶`: [u8(0xE5), 0xB8] // U+87F6 <cjk>
	`蟷`: [u8(0xE5), 0xB9] // U+87F7 <cjk>
	`蠎`: [u8(0xE5), 0xBA] // U+880E <cjk>
	`蟒`: [u8(0xE5), 0xBB] // U+87D2 <cjk>
	`蠑`: [u8(0xE5), 0xBC] // U+8811 <cjk>
	`蠖`: [u8(0xE5), 0xBD] // U+8816 <cjk>
	`蠕`: [u8(0xE5), 0xBE] // U+8815 <cjk>
	`蠢`: [u8(0xE5), 0xBF] // U+8822 <cjk>
	`蠡`: [u8(0xE5), 0xC0] // U+8821 <cjk>
	`蠱`: [u8(0xE5), 0xC1] // U+8831 <cjk>
	`蠶`: [u8(0xE5), 0xC2] // U+8836 <cjk>
	`蠹`: [u8(0xE5), 0xC3] // U+8839 <cjk>
	`蠧`: [u8(0xE5), 0xC4] // U+8827 <cjk>
	`蠻`: [u8(0xE5), 0xC5] // U+883B <cjk>
	`衄`: [u8(0xE5), 0xC6] // U+8844 <cjk>
	`衂`: [u8(0xE5), 0xC7] // U+8842 <cjk>
	`衒`: [u8(0xE5), 0xC8] // U+8852 <cjk>
	`衙`: [u8(0xE5), 0xC9] // U+8859 <cjk>
	`衞`: [u8(0xE5), 0xCA] // U+885E <cjk>
	`衢`: [u8(0xE5), 0xCB] // U+8862 <cjk>
	`衫`: [u8(0xE5), 0xCC] // U+886B <cjk>
	`袁`: [u8(0xE5), 0xCD] // U+8881 <cjk>
	`衾`: [u8(0xE5), 0xCE] // U+887E <cjk>
	`袞`: [u8(0xE5), 0xCF] // U+889E <cjk>
	`衵`: [u8(0xE5), 0xD0] // U+8875 <cjk>
	`衽`: [u8(0xE5), 0xD1] // U+887D <cjk>
	`袵`: [u8(0xE5), 0xD2] // U+88B5 <cjk>
	`衲`: [u8(0xE5), 0xD3] // U+8872 <cjk>
	`袂`: [u8(0xE5), 0xD4] // U+8882 <cjk>
	`袗`: [u8(0xE5), 0xD5] // U+8897 <cjk>
	`袒`: [u8(0xE5), 0xD6] // U+8892 <cjk>
	`袮`: [u8(0xE5), 0xD7] // U+88AE <cjk>
	`袙`: [u8(0xE5), 0xD8] // U+8899 <cjk>
	`袢`: [u8(0xE5), 0xD9] // U+88A2 <cjk>
	`袍`: [u8(0xE5), 0xDA] // U+888D <cjk>
	`袤`: [u8(0xE5), 0xDB] // U+88A4 <cjk>
	`袰`: [u8(0xE5), 0xDC] // U+88B0 <cjk>
	`袿`: [u8(0xE5), 0xDD] // U+88BF <cjk>
	`袱`: [u8(0xE5), 0xDE] // U+88B1 <cjk>
	`裃`: [u8(0xE5), 0xDF] // U+88C3 <cjk>
	`裄`: [u8(0xE5), 0xE0] // U+88C4 <cjk>
	`裔`: [u8(0xE5), 0xE1] // U+88D4 <cjk>
	`裘`: [u8(0xE5), 0xE2] // U+88D8 <cjk>
	`裙`: [u8(0xE5), 0xE3] // U+88D9 <cjk>
	`裝`: [u8(0xE5), 0xE4] // U+88DD <cjk>
	`裹`: [u8(0xE5), 0xE5] // U+88F9 <cjk>
	`褂`: [u8(0xE5), 0xE6] // U+8902 <cjk>
	`裼`: [u8(0xE5), 0xE7] // U+88FC <cjk>
	`裴`: [u8(0xE5), 0xE8] // U+88F4 <cjk>
	`裨`: [u8(0xE5), 0xE9] // U+88E8 <cjk>
	`裲`: [u8(0xE5), 0xEA] // U+88F2 <cjk>
	`褄`: [u8(0xE5), 0xEB] // U+8904 <cjk>
	`褌`: [u8(0xE5), 0xEC] // U+890C <cjk>
	`褊`: [u8(0xE5), 0xED] // U+890A <cjk>
	`褓`: [u8(0xE5), 0xEE] // U+8913 <cjk>
	`襃`: [u8(0xE5), 0xEF] // U+8943 <cjk>
	`褞`: [u8(0xE5), 0xF0] // U+891E <cjk>
	`褥`: [u8(0xE5), 0xF1] // U+8925 <cjk>
	`褪`: [u8(0xE5), 0xF2] // U+892A <cjk>
	`褫`: [u8(0xE5), 0xF3] // U+892B <cjk>
	`襁`: [u8(0xE5), 0xF4] // U+8941 <cjk>
	`襄`: [u8(0xE5), 0xF5] // U+8944 <cjk>
	`褻`: [u8(0xE5), 0xF6] // U+893B <cjk>
	`褶`: [u8(0xE5), 0xF7] // U+8936 <cjk>
	`褸`: [u8(0xE5), 0xF8] // U+8938 <cjk>
	`襌`: [u8(0xE5), 0xF9] // U+894C <cjk>
	`褝`: [u8(0xE5), 0xFA] // U+891D <cjk>
	`襠`: [u8(0xE5), 0xFB] // U+8960 <cjk>
	`襞`: [u8(0xE5), 0xFC] // U+895E <cjk>
	`襦`: [u8(0xE6), 0x40] // U+8966 <cjk>
	`襤`: [u8(0xE6), 0x41] // U+8964 <cjk>
	`襭`: [u8(0xE6), 0x42] // U+896D <cjk>
	`襪`: [u8(0xE6), 0x43] // U+896A <cjk>
	`襯`: [u8(0xE6), 0x44] // U+896F <cjk>
	`襴`: [u8(0xE6), 0x45] // U+8974 <cjk>
	`襷`: [u8(0xE6), 0x46] // U+8977 <cjk>
	`襾`: [u8(0xE6), 0x47] // U+897E <cjk>
	`覃`: [u8(0xE6), 0x48] // U+8983 <cjk>
	`覈`: [u8(0xE6), 0x49] // U+8988 <cjk>
	`覊`: [u8(0xE6), 0x4A] // U+898A <cjk>
	`覓`: [u8(0xE6), 0x4B] // U+8993 <cjk>
	`覘`: [u8(0xE6), 0x4C] // U+8998 <cjk>
	`覡`: [u8(0xE6), 0x4D] // U+89A1 <cjk>
	`覩`: [u8(0xE6), 0x4E] // U+89A9 <cjk>
	`覦`: [u8(0xE6), 0x4F] // U+89A6 <cjk>
	`覬`: [u8(0xE6), 0x50] // U+89AC <cjk>
	`覯`: [u8(0xE6), 0x51] // U+89AF <cjk>
	`覲`: [u8(0xE6), 0x52] // U+89B2 <cjk>
	`覺`: [u8(0xE6), 0x53] // U+89BA <cjk>
	`覽`: [u8(0xE6), 0x54] // U+89BD <cjk>
	`覿`: [u8(0xE6), 0x55] // U+89BF <cjk>
	`觀`: [u8(0xE6), 0x56] // U+89C0 <cjk>
	`觚`: [u8(0xE6), 0x57] // U+89DA <cjk>
	`觜`: [u8(0xE6), 0x58] // U+89DC <cjk>
	`觝`: [u8(0xE6), 0x59] // U+89DD <cjk>
	`觧`: [u8(0xE6), 0x5A] // U+89E7 <cjk>
	`觴`: [u8(0xE6), 0x5B] // U+89F4 <cjk>
	`觸`: [u8(0xE6), 0x5C] // U+89F8 <cjk>
	`訃`: [u8(0xE6), 0x5D] // U+8A03 <cjk>
	`訖`: [u8(0xE6), 0x5E] // U+8A16 <cjk>
	`訐`: [u8(0xE6), 0x5F] // U+8A10 <cjk>
	`訌`: [u8(0xE6), 0x60] // U+8A0C <cjk>
	`訛`: [u8(0xE6), 0x61] // U+8A1B <cjk>
	`訝`: [u8(0xE6), 0x62] // U+8A1D <cjk>
	`訥`: [u8(0xE6), 0x63] // U+8A25 <cjk>
	`訶`: [u8(0xE6), 0x64] // U+8A36 <cjk>
	`詁`: [u8(0xE6), 0x65] // U+8A41 <cjk>
	`詛`: [u8(0xE6), 0x66] // U+8A5B <cjk>
	`詒`: [u8(0xE6), 0x67] // U+8A52 <cjk>
	`詆`: [u8(0xE6), 0x68] // U+8A46 <cjk>
	`詈`: [u8(0xE6), 0x69] // U+8A48 <cjk>
	`詼`: [u8(0xE6), 0x6A] // U+8A7C <cjk>
	`詭`: [u8(0xE6), 0x6B] // U+8A6D <cjk>
	`詬`: [u8(0xE6), 0x6C] // U+8A6C <cjk>
	`詢`: [u8(0xE6), 0x6D] // U+8A62 <cjk>
	`誅`: [u8(0xE6), 0x6E] // U+8A85 <cjk>
	`誂`: [u8(0xE6), 0x6F] // U+8A82 <cjk>
	`誄`: [u8(0xE6), 0x70] // U+8A84 <cjk>
	`誨`: [u8(0xE6), 0x71] // U+8AA8 <cjk>
	`誡`: [u8(0xE6), 0x72] // U+8AA1 <cjk>
	`誑`: [u8(0xE6), 0x73] // U+8A91 <cjk>
	`誥`: [u8(0xE6), 0x74] // U+8AA5 <cjk>
	`誦`: [u8(0xE6), 0x75] // U+8AA6 <cjk>
	`誚`: [u8(0xE6), 0x76] // U+8A9A <cjk>
	`誣`: [u8(0xE6), 0x77] // U+8AA3 <cjk>
	`諄`: [u8(0xE6), 0x78] // U+8AC4 <cjk>
	`諍`: [u8(0xE6), 0x79] // U+8ACD <cjk>
	`諂`: [u8(0xE6), 0x7A] // U+8AC2 <cjk>
	`諚`: [u8(0xE6), 0x7B] // U+8ADA <cjk>
	`諫`: [u8(0xE6), 0x7C] // U+8AEB <cjk>
	`諳`: [u8(0xE6), 0x7D] // U+8AF3 <cjk>
	`諧`: [u8(0xE6), 0x7E] // U+8AE7 <cjk>
	`諤`: [u8(0xE6), 0x80] // U+8AE4 <cjk>
	`諱`: [u8(0xE6), 0x81] // U+8AF1 <cjk>
	`謔`: [u8(0xE6), 0x82] // U+8B14 <cjk>
	`諠`: [u8(0xE6), 0x83] // U+8AE0 <cjk>
	`諢`: [u8(0xE6), 0x84] // U+8AE2 <cjk>
	`諷`: [u8(0xE6), 0x85] // U+8AF7 <cjk>
	`諞`: [u8(0xE6), 0x86] // U+8ADE <cjk>
	`諛`: [u8(0xE6), 0x87] // U+8ADB <cjk>
	`謌`: [u8(0xE6), 0x88] // U+8B0C <cjk>
	`謇`: [u8(0xE6), 0x89] // U+8B07 <cjk>
	`謚`: [u8(0xE6), 0x8A] // U+8B1A <cjk>
	`諡`: [u8(0xE6), 0x8B] // U+8AE1 <cjk>
	`謖`: [u8(0xE6), 0x8C] // U+8B16 <cjk>
	`謐`: [u8(0xE6), 0x8D] // U+8B10 <cjk>
	`謗`: [u8(0xE6), 0x8E] // U+8B17 <cjk>
	`謠`: [u8(0xE6), 0x8F] // U+8B20 <cjk>
	`謳`: [u8(0xE6), 0x90] // U+8B33 <cjk>
	`鞫`: [u8(0xE6), 0x91] // U+97AB <cjk>
	`謦`: [u8(0xE6), 0x92] // U+8B26 <cjk>
	`謫`: [u8(0xE6), 0x93] // U+8B2B <cjk>
	`謾`: [u8(0xE6), 0x94] // U+8B3E <cjk>
	`謨`: [u8(0xE6), 0x95] // U+8B28 <cjk>
	`譁`: [u8(0xE6), 0x96] // U+8B41 <cjk>
	`譌`: [u8(0xE6), 0x97] // U+8B4C <cjk>
	`譏`: [u8(0xE6), 0x98] // U+8B4F <cjk>
	`譎`: [u8(0xE6), 0x99] // U+8B4E <cjk>
	`證`: [u8(0xE6), 0x9A] // U+8B49 <cjk>
	`譖`: [u8(0xE6), 0x9B] // U+8B56 <cjk>
	`譛`: [u8(0xE6), 0x9C] // U+8B5B <cjk>
	`譚`: [u8(0xE6), 0x9D] // U+8B5A <cjk>
	`譫`: [u8(0xE6), 0x9E] // U+8B6B <cjk>
	`譟`: [u8(0xE6), 0x9F] // U+8B5F <cjk>
	`譬`: [u8(0xE6), 0xA0] // U+8B6C <cjk>
	`譯`: [u8(0xE6), 0xA1] // U+8B6F <cjk>
	`譴`: [u8(0xE6), 0xA2] // U+8B74 <cjk>
	`譽`: [u8(0xE6), 0xA3] // U+8B7D <cjk>
	`讀`: [u8(0xE6), 0xA4] // U+8B80 <cjk>
	`讌`: [u8(0xE6), 0xA5] // U+8B8C <cjk>
	`讎`: [u8(0xE6), 0xA6] // U+8B8E <cjk>
	`讒`: [u8(0xE6), 0xA7] // U+8B92 <cjk>
	`讓`: [u8(0xE6), 0xA8] // U+8B93 <cjk>
	`讖`: [u8(0xE6), 0xA9] // U+8B96 <cjk>
	`讙`: [u8(0xE6), 0xAA] // U+8B99 <cjk>
	`讚`: [u8(0xE6), 0xAB] // U+8B9A <cjk>
	`谺`: [u8(0xE6), 0xAC] // U+8C3A <cjk>
	`豁`: [u8(0xE6), 0xAD] // U+8C41 <cjk>
	`谿`: [u8(0xE6), 0xAE] // U+8C3F <cjk>
	`豈`: [u8(0xE6), 0xAF] // U+8C48 <cjk>
	`豌`: [u8(0xE6), 0xB0] // U+8C4C <cjk>
	`豎`: [u8(0xE6), 0xB1] // U+8C4E <cjk>
	`豐`: [u8(0xE6), 0xB2] // U+8C50 <cjk>
	`豕`: [u8(0xE6), 0xB3] // U+8C55 <cjk>
	`豢`: [u8(0xE6), 0xB4] // U+8C62 <cjk>
	`豬`: [u8(0xE6), 0xB5] // U+8C6C <cjk>
	`豸`: [u8(0xE6), 0xB6] // U+8C78 <cjk>
	`豺`: [u8(0xE6), 0xB7] // U+8C7A <cjk>
	`貂`: [u8(0xE6), 0xB8] // U+8C82 <cjk>
	`貉`: [u8(0xE6), 0xB9] // U+8C89 <cjk>
	`貅`: [u8(0xE6), 0xBA] // U+8C85 <cjk>
	`貊`: [u8(0xE6), 0xBB] // U+8C8A <cjk>
	`貍`: [u8(0xE6), 0xBC] // U+8C8D <cjk>
	`貎`: [u8(0xE6), 0xBD] // U+8C8E <cjk>
	`貔`: [u8(0xE6), 0xBE] // U+8C94 <cjk>
	`豼`: [u8(0xE6), 0xBF] // U+8C7C <cjk>
	`貘`: [u8(0xE6), 0xC0] // U+8C98 <cjk>
	`戝`: [u8(0xE6), 0xC1] // U+621D <cjk>
	`貭`: [u8(0xE6), 0xC2] // U+8CAD <cjk>
	`貪`: [u8(0xE6), 0xC3] // U+8CAA <cjk>
	`貽`: [u8(0xE6), 0xC4] // U+8CBD <cjk>
	`貲`: [u8(0xE6), 0xC5] // U+8CB2 <cjk>
	`貳`: [u8(0xE6), 0xC6] // U+8CB3 <cjk>
	`貮`: [u8(0xE6), 0xC7] // U+8CAE <cjk>
	`貶`: [u8(0xE6), 0xC8] // U+8CB6 <cjk>
	`賈`: [u8(0xE6), 0xC9] // U+8CC8 <cjk>
	`賁`: [u8(0xE6), 0xCA] // U+8CC1 <cjk>
	`賤`: [u8(0xE6), 0xCB] // U+8CE4 <cjk>
	`賣`: [u8(0xE6), 0xCC] // U+8CE3 <cjk>
	`賚`: [u8(0xE6), 0xCD] // U+8CDA <cjk>
	`賽`: [u8(0xE6), 0xCE] // U+8CFD <cjk>
	`賺`: [u8(0xE6), 0xCF] // U+8CFA <cjk>
	`賻`: [u8(0xE6), 0xD0] // U+8CFB <cjk>
	`贄`: [u8(0xE6), 0xD1] // U+8D04 <cjk>
	`贅`: [u8(0xE6), 0xD2] // U+8D05 <cjk>
	`贊`: [u8(0xE6), 0xD3] // U+8D0A <cjk>
	`贇`: [u8(0xE6), 0xD4] // U+8D07 <cjk>
	`贏`: [u8(0xE6), 0xD5] // U+8D0F <cjk>
	`贍`: [u8(0xE6), 0xD6] // U+8D0D <cjk>
	`贐`: [u8(0xE6), 0xD7] // U+8D10 <cjk>
	`齎`: [u8(0xE6), 0xD8] // U+9F4E <cjk>
	`贓`: [u8(0xE6), 0xD9] // U+8D13 <cjk>
	`賍`: [u8(0xE6), 0xDA] // U+8CCD <cjk>
	`贔`: [u8(0xE6), 0xDB] // U+8D14 <cjk>
	`贖`: [u8(0xE6), 0xDC] // U+8D16 <cjk>
	`赧`: [u8(0xE6), 0xDD] // U+8D67 <cjk>
	`赭`: [u8(0xE6), 0xDE] // U+8D6D <cjk>
	`赱`: [u8(0xE6), 0xDF] // U+8D71 <cjk>
	`赳`: [u8(0xE6), 0xE0] // U+8D73 <cjk>
	`趁`: [u8(0xE6), 0xE1] // U+8D81 <cjk>
	`趙`: [u8(0xE6), 0xE2] // U+8D99 <cjk>
	`跂`: [u8(0xE6), 0xE3] // U+8DC2 <cjk>
	`趾`: [u8(0xE6), 0xE4] // U+8DBE <cjk>
	`趺`: [u8(0xE6), 0xE5] // U+8DBA <cjk>
	`跏`: [u8(0xE6), 0xE6] // U+8DCF <cjk>
	`跚`: [u8(0xE6), 0xE7] // U+8DDA <cjk>
	`跖`: [u8(0xE6), 0xE8] // U+8DD6 <cjk>
	`跌`: [u8(0xE6), 0xE9] // U+8DCC <cjk>
	`跛`: [u8(0xE6), 0xEA] // U+8DDB <cjk>
	`跋`: [u8(0xE6), 0xEB] // U+8DCB <cjk>
	`跪`: [u8(0xE6), 0xEC] // U+8DEA <cjk>
	`跫`: [u8(0xE6), 0xED] // U+8DEB <cjk>
	`跟`: [u8(0xE6), 0xEE] // U+8DDF <cjk>
	`跣`: [u8(0xE6), 0xEF] // U+8DE3 <cjk>
	`跼`: [u8(0xE6), 0xF0] // U+8DFC <cjk>
	`踈`: [u8(0xE6), 0xF1] // U+8E08 <cjk>
	`踉`: [u8(0xE6), 0xF2] // U+8E09 <cjk>
	`跿`: [u8(0xE6), 0xF3] // U+8DFF <cjk>
	`踝`: [u8(0xE6), 0xF4] // U+8E1D <cjk>
	`踞`: [u8(0xE6), 0xF5] // U+8E1E <cjk>
	`踐`: [u8(0xE6), 0xF6] // U+8E10 <cjk>
	`踟`: [u8(0xE6), 0xF7] // U+8E1F <cjk>
	`蹂`: [u8(0xE6), 0xF8] // U+8E42 <cjk>
	`踵`: [u8(0xE6), 0xF9] // U+8E35 <cjk>
	`踰`: [u8(0xE6), 0xFA] // U+8E30 <cjk>
	`踴`: [u8(0xE6), 0xFB] // U+8E34 <cjk>
	`蹊`: [u8(0xE6), 0xFC] // U+8E4A <cjk>
	`蹇`: [u8(0xE7), 0x40] // U+8E47 <cjk>
	`蹉`: [u8(0xE7), 0x41] // U+8E49 <cjk>
	`蹌`: [u8(0xE7), 0x42] // U+8E4C <cjk>
	`蹐`: [u8(0xE7), 0x43] // U+8E50 <cjk>
	`蹈`: [u8(0xE7), 0x44] // U+8E48 <cjk>
	`蹙`: [u8(0xE7), 0x45] // U+8E59 <cjk>
	`蹤`: [u8(0xE7), 0x46] // U+8E64 <cjk>
	`蹠`: [u8(0xE7), 0x47] // U+8E60 <cjk>
	`踪`: [u8(0xE7), 0x48] // U+8E2A <cjk>
	`蹣`: [u8(0xE7), 0x49] // U+8E63 <cjk>
	`蹕`: [u8(0xE7), 0x4A] // U+8E55 <cjk>
	`蹶`: [u8(0xE7), 0x4B] // U+8E76 <cjk>
	`蹲`: [u8(0xE7), 0x4C] // U+8E72 <cjk>
	`蹼`: [u8(0xE7), 0x4D] // U+8E7C <cjk>
	`躁`: [u8(0xE7), 0x4E] // U+8E81 <cjk>
	`躇`: [u8(0xE7), 0x4F] // U+8E87 <cjk>
	`躅`: [u8(0xE7), 0x50] // U+8E85 <cjk>
	`躄`: [u8(0xE7), 0x51] // U+8E84 <cjk>
	`躋`: [u8(0xE7), 0x52] // U+8E8B <cjk>
	`躊`: [u8(0xE7), 0x53] // U+8E8A <cjk>
	`躓`: [u8(0xE7), 0x54] // U+8E93 <cjk>
	`躑`: [u8(0xE7), 0x55] // U+8E91 <cjk>
	`躔`: [u8(0xE7), 0x56] // U+8E94 <cjk>
	`躙`: [u8(0xE7), 0x57] // U+8E99 <cjk>
	`躪`: [u8(0xE7), 0x58] // U+8EAA <cjk>
	`躡`: [u8(0xE7), 0x59] // U+8EA1 <cjk>
	`躬`: [u8(0xE7), 0x5A] // U+8EAC <cjk>
	`躰`: [u8(0xE7), 0x5B] // U+8EB0 <cjk>
	`軆`: [u8(0xE7), 0x5C] // U+8EC6 <cjk>
	`躱`: [u8(0xE7), 0x5D] // U+8EB1 <cjk>
	`躾`: [u8(0xE7), 0x5E] // U+8EBE <cjk>
	`軅`: [u8(0xE7), 0x5F] // U+8EC5 <cjk>
	`軈`: [u8(0xE7), 0x60] // U+8EC8 <cjk>
	`軋`: [u8(0xE7), 0x61] // U+8ECB <cjk>
	`軛`: [u8(0xE7), 0x62] // U+8EDB <cjk>
	`軣`: [u8(0xE7), 0x63] // U+8EE3 <cjk>
	`軼`: [u8(0xE7), 0x64] // U+8EFC <cjk>
	`軻`: [u8(0xE7), 0x65] // U+8EFB <cjk>
	`軫`: [u8(0xE7), 0x66] // U+8EEB <cjk>
	`軾`: [u8(0xE7), 0x67] // U+8EFE <cjk>
	`輊`: [u8(0xE7), 0x68] // U+8F0A <cjk>
	`輅`: [u8(0xE7), 0x69] // U+8F05 <cjk>
	`輕`: [u8(0xE7), 0x6A] // U+8F15 <cjk>
	`輒`: [u8(0xE7), 0x6B] // U+8F12 <cjk>
	`輙`: [u8(0xE7), 0x6C] // U+8F19 <cjk>
	`輓`: [u8(0xE7), 0x6D] // U+8F13 <cjk>
	`輜`: [u8(0xE7), 0x6E] // U+8F1C <cjk>
	`輟`: [u8(0xE7), 0x6F] // U+8F1F <cjk>
	`輛`: [u8(0xE7), 0x70] // U+8F1B <cjk>
	`輌`: [u8(0xE7), 0x71] // U+8F0C <cjk>
	`輦`: [u8(0xE7), 0x72] // U+8F26 <cjk>
	`輳`: [u8(0xE7), 0x73] // U+8F33 <cjk>
	`輻`: [u8(0xE7), 0x74] // U+8F3B <cjk>
	`輹`: [u8(0xE7), 0x75] // U+8F39 <cjk>
	`轅`: [u8(0xE7), 0x76] // U+8F45 <cjk>
	`轂`: [u8(0xE7), 0x77] // U+8F42 <cjk>
	`輾`: [u8(0xE7), 0x78] // U+8F3E <cjk>
	`轌`: [u8(0xE7), 0x79] // U+8F4C <cjk>
	`轉`: [u8(0xE7), 0x7A] // U+8F49 <cjk>
	`轆`: [u8(0xE7), 0x7B] // U+8F46 <cjk>
	`轎`: [u8(0xE7), 0x7C] // U+8F4E <cjk>
	`轗`: [u8(0xE7), 0x7D] // U+8F57 <cjk>
	`轜`: [u8(0xE7), 0x7E] // U+8F5C <cjk>
	`轢`: [u8(0xE7), 0x80] // U+8F62 <cjk>
	`轣`: [u8(0xE7), 0x81] // U+8F63 <cjk>
	`轤`: [u8(0xE7), 0x82] // U+8F64 <cjk>
	`辜`: [u8(0xE7), 0x83] // U+8F9C <cjk>
	`辟`: [u8(0xE7), 0x84] // U+8F9F <cjk>
	`辣`: [u8(0xE7), 0x85] // U+8FA3 <cjk>
	`辭`: [u8(0xE7), 0x86] // U+8FAD <cjk>
	`辯`: [u8(0xE7), 0x87] // U+8FAF <cjk>
	`辷`: [u8(0xE7), 0x88] // U+8FB7 <cjk>
	`迚`: [u8(0xE7), 0x89] // U+8FDA <cjk>
	`迥`: [u8(0xE7), 0x8A] // U+8FE5 <cjk>
	`迢`: [u8(0xE7), 0x8B] // U+8FE2 <cjk>
	`迪`: [u8(0xE7), 0x8C] // U+8FEA <cjk>
	`迯`: [u8(0xE7), 0x8D] // U+8FEF <cjk>
	`邇`: [u8(0xE7), 0x8E] // U+9087 <cjk>
	`迴`: [u8(0xE7), 0x8F] // U+8FF4 <cjk>
	`逅`: [u8(0xE7), 0x90] // U+9005 <cjk>
	`迹`: [u8(0xE7), 0x91] // U+8FF9 <cjk>
	`迺`: [u8(0xE7), 0x92] // U+8FFA <cjk>
	`逑`: [u8(0xE7), 0x93] // U+9011 <cjk>
	`逕`: [u8(0xE7), 0x94] // U+9015 <cjk>
	`逡`: [u8(0xE7), 0x95] // U+9021 <cjk>
	`逍`: [u8(0xE7), 0x96] // U+900D <cjk>
	`逞`: [u8(0xE7), 0x97] // U+901E <cjk>
	`逖`: [u8(0xE7), 0x98] // U+9016 <cjk>
	`逋`: [u8(0xE7), 0x99] // U+900B <cjk>
	`逧`: [u8(0xE7), 0x9A] // U+9027 <cjk>
	`逶`: [u8(0xE7), 0x9B] // U+9036 <cjk>
	`逵`: [u8(0xE7), 0x9C] // U+9035 <cjk>
	`逹`: [u8(0xE7), 0x9D] // U+9039 <cjk>
	`迸`: [u8(0xE7), 0x9E] // U+8FF8 <cjk>
	`遏`: [u8(0xE7), 0x9F] // U+904F <cjk>
	`遐`: [u8(0xE7), 0xA0] // U+9050 <cjk>
	`遑`: [u8(0xE7), 0xA1] // U+9051 <cjk>
	`遒`: [u8(0xE7), 0xA2] // U+9052 <cjk>
	`逎`: [u8(0xE7), 0xA3] // U+900E <cjk>
	`遉`: [u8(0xE7), 0xA4] // U+9049 <cjk>
	`逾`: [u8(0xE7), 0xA5] // U+903E <cjk>
	`遖`: [u8(0xE7), 0xA6] // U+9056 <cjk>
	`遘`: [u8(0xE7), 0xA7] // U+9058 <cjk>
	`遞`: [u8(0xE7), 0xA8] // U+905E <cjk>
	`遨`: [u8(0xE7), 0xA9] // U+9068 <cjk>
	`遯`: [u8(0xE7), 0xAA] // U+906F <cjk>
	`遶`: [u8(0xE7), 0xAB] // U+9076 <cjk>
	`隨`: [u8(0xE7), 0xAC] // U+96A8 <cjk>
	`遲`: [u8(0xE7), 0xAD] // U+9072 <cjk>
	`邂`: [u8(0xE7), 0xAE] // U+9082 <cjk>
	`遽`: [u8(0xE7), 0xAF] // U+907D <cjk>
	`邁`: [u8(0xE7), 0xB0] // U+9081 <cjk>
	`邀`: [u8(0xE7), 0xB1] // U+9080 <cjk>
	`邊`: [u8(0xE7), 0xB2] // U+908A <cjk>
	`邉`: [u8(0xE7), 0xB3] // U+9089 <cjk>
	`邏`: [u8(0xE7), 0xB4] // U+908F <cjk>
	`邨`: [u8(0xE7), 0xB5] // U+90A8 <cjk>
	`邯`: [u8(0xE7), 0xB6] // U+90AF <cjk>
	`邱`: [u8(0xE7), 0xB7] // U+90B1 <cjk>
	`邵`: [u8(0xE7), 0xB8] // U+90B5 <cjk>
	`郢`: [u8(0xE7), 0xB9] // U+90E2 <cjk>
	`郤`: [u8(0xE7), 0xBA] // U+90E4 <cjk>
	`扈`: [u8(0xE7), 0xBB] // U+6248 <cjk>
	`郛`: [u8(0xE7), 0xBC] // U+90DB <cjk>
	`鄂`: [u8(0xE7), 0xBD] // U+9102 <cjk>
	`鄒`: [u8(0xE7), 0xBE] // U+9112 <cjk>
	`鄙`: [u8(0xE7), 0xBF] // U+9119 <cjk>
	`鄲`: [u8(0xE7), 0xC0] // U+9132 <cjk>
	`鄰`: [u8(0xE7), 0xC1] // U+9130 <cjk>
	`酊`: [u8(0xE7), 0xC2] // U+914A <cjk>
	`酖`: [u8(0xE7), 0xC3] // U+9156 <cjk>
	`酘`: [u8(0xE7), 0xC4] // U+9158 <cjk>
	`酣`: [u8(0xE7), 0xC5] // U+9163 <cjk>
	`酥`: [u8(0xE7), 0xC6] // U+9165 <cjk>
	`酩`: [u8(0xE7), 0xC7] // U+9169 <cjk>
	`酳`: [u8(0xE7), 0xC8] // U+9173 <cjk>
	`酲`: [u8(0xE7), 0xC9] // U+9172 <cjk>
	`醋`: [u8(0xE7), 0xCA] // U+918B <cjk>
	`醉`: [u8(0xE7), 0xCB] // U+9189 <cjk>
	`醂`: [u8(0xE7), 0xCC] // U+9182 <cjk>
	`醢`: [u8(0xE7), 0xCD] // U+91A2 <cjk>
	`醫`: [u8(0xE7), 0xCE] // U+91AB <cjk>
	`醯`: [u8(0xE7), 0xCF] // U+91AF <cjk>
	`醪`: [u8(0xE7), 0xD0] // U+91AA <cjk>
	`醵`: [u8(0xE7), 0xD1] // U+91B5 <cjk>
	`醴`: [u8(0xE7), 0xD2] // U+91B4 <cjk>
	`醺`: [u8(0xE7), 0xD3] // U+91BA <cjk>
	`釀`: [u8(0xE7), 0xD4] // U+91C0 <cjk>
	`釁`: [u8(0xE7), 0xD5] // U+91C1 <cjk>
	`釉`: [u8(0xE7), 0xD6] // U+91C9 <cjk>
	`釋`: [u8(0xE7), 0xD7] // U+91CB <cjk>
	`釐`: [u8(0xE7), 0xD8] // U+91D0 <cjk>
	`釖`: [u8(0xE7), 0xD9] // U+91D6 <cjk>
	`釟`: [u8(0xE7), 0xDA] // U+91DF <cjk>
	`釡`: [u8(0xE7), 0xDB] // U+91E1 <cjk>
	`釛`: [u8(0xE7), 0xDC] // U+91DB <cjk>
	`釼`: [u8(0xE7), 0xDD] // U+91FC <cjk>
	`釵`: [u8(0xE7), 0xDE] // U+91F5 <cjk>
	`釶`: [u8(0xE7), 0xDF] // U+91F6 <cjk>
	`鈞`: [u8(0xE7), 0xE0] // U+921E <cjk>
	`釿`: [u8(0xE7), 0xE1] // U+91FF <cjk>
	`鈔`: [u8(0xE7), 0xE2] // U+9214 <cjk>
	`鈬`: [u8(0xE7), 0xE3] // U+922C <cjk>
	`鈕`: [u8(0xE7), 0xE4] // U+9215 <cjk>
	`鈑`: [u8(0xE7), 0xE5] // U+9211 <cjk>
	`鉞`: [u8(0xE7), 0xE6] // U+925E <cjk>
	`鉗`: [u8(0xE7), 0xE7] // U+9257 <cjk>
	`鉅`: [u8(0xE7), 0xE8] // U+9245 <cjk>
	`鉉`: [u8(0xE7), 0xE9] // U+9249 <cjk>
	`鉤`: [u8(0xE7), 0xEA] // U+9264 <cjk>
	`鉈`: [u8(0xE7), 0xEB] // U+9248 <cjk>
	`銕`: [u8(0xE7), 0xEC] // U+9295 <cjk>
	`鈿`: [u8(0xE7), 0xED] // U+923F <cjk>
	`鉋`: [u8(0xE7), 0xEE] // U+924B <cjk>
	`鉐`: [u8(0xE7), 0xEF] // U+9250 <cjk>
	`銜`: [u8(0xE7), 0xF0] // U+929C <cjk>
	`銖`: [u8(0xE7), 0xF1] // U+9296 <cjk>
	`銓`: [u8(0xE7), 0xF2] // U+9293 <cjk>
	`銛`: [u8(0xE7), 0xF3] // U+929B <cjk>
	`鉚`: [u8(0xE7), 0xF4] // U+925A <cjk>
	`鋏`: [u8(0xE7), 0xF5] // U+92CF <cjk>
	`銹`: [u8(0xE7), 0xF6] // U+92B9 <cjk>
	`銷`: [u8(0xE7), 0xF7] // U+92B7 <cjk>
	`鋩`: [u8(0xE7), 0xF8] // U+92E9 <cjk>
	`錏`: [u8(0xE7), 0xF9] // U+930F <cjk>
	`鋺`: [u8(0xE7), 0xFA] // U+92FA <cjk>
	`鍄`: [u8(0xE7), 0xFB] // U+9344 <cjk>
	`錮`: [u8(0xE7), 0xFC] // U+932E <cjk>
	`錙`: [u8(0xE8), 0x40] // U+9319 <cjk>
	`錢`: [u8(0xE8), 0x41] // U+9322 <cjk>
	`錚`: [u8(0xE8), 0x42] // U+931A <cjk>
	`錣`: [u8(0xE8), 0x43] // U+9323 <cjk>
	`錺`: [u8(0xE8), 0x44] // U+933A <cjk>
	`錵`: [u8(0xE8), 0x45] // U+9335 <cjk>
	`錻`: [u8(0xE8), 0x46] // U+933B <cjk>
	`鍜`: [u8(0xE8), 0x47] // U+935C <cjk>
	`鍠`: [u8(0xE8), 0x48] // U+9360 <cjk>
	`鍼`: [u8(0xE8), 0x49] // U+937C <cjk>
	`鍮`: [u8(0xE8), 0x4A] // U+936E <cjk>
	`鍖`: [u8(0xE8), 0x4B] // U+9356 <cjk>
	`鎰`: [u8(0xE8), 0x4C] // U+93B0 <cjk>
	`鎬`: [u8(0xE8), 0x4D] // U+93AC <cjk>
	`鎭`: [u8(0xE8), 0x4E] // U+93AD <cjk>
	`鎔`: [u8(0xE8), 0x4F] // U+9394 <cjk>
	`鎹`: [u8(0xE8), 0x50] // U+93B9 <cjk>
	`鏖`: [u8(0xE8), 0x51] // U+93D6 <cjk>
	`鏗`: [u8(0xE8), 0x52] // U+93D7 <cjk>
	`鏨`: [u8(0xE8), 0x53] // U+93E8 <cjk>
	`鏥`: [u8(0xE8), 0x54] // U+93E5 <cjk>
	`鏘`: [u8(0xE8), 0x55] // U+93D8 <cjk>
	`鏃`: [u8(0xE8), 0x56] // U+93C3 <cjk>
	`鏝`: [u8(0xE8), 0x57] // U+93DD <cjk>
	`鏐`: [u8(0xE8), 0x58] // U+93D0 <cjk>
	`鏈`: [u8(0xE8), 0x59] // U+93C8 <cjk>
	`鏤`: [u8(0xE8), 0x5A] // U+93E4 <cjk>
	`鐚`: [u8(0xE8), 0x5B] // U+941A <cjk>
	`鐔`: [u8(0xE8), 0x5C] // U+9414 <cjk>
	`鐓`: [u8(0xE8), 0x5D] // U+9413 <cjk>
	`鐃`: [u8(0xE8), 0x5E] // U+9403 <cjk>
	`鐇`: [u8(0xE8), 0x5F] // U+9407 <cjk>
	`鐐`: [u8(0xE8), 0x60] // U+9410 <cjk>
	`鐶`: [u8(0xE8), 0x61] // U+9436 <cjk>
	`鐫`: [u8(0xE8), 0x62] // U+942B <cjk>
	`鐵`: [u8(0xE8), 0x63] // U+9435 <cjk>
	`鐡`: [u8(0xE8), 0x64] // U+9421 <cjk>
	`鐺`: [u8(0xE8), 0x65] // U+943A <cjk>
	`鑁`: [u8(0xE8), 0x66] // U+9441 <cjk>
	`鑒`: [u8(0xE8), 0x67] // U+9452 <cjk>
	`鑄`: [u8(0xE8), 0x68] // U+9444 <cjk>
	`鑛`: [u8(0xE8), 0x69] // U+945B <cjk>
	`鑠`: [u8(0xE8), 0x6A] // U+9460 <cjk>
	`鑢`: [u8(0xE8), 0x6B] // U+9462 <cjk>
	`鑞`: [u8(0xE8), 0x6C] // U+945E <cjk>
	`鑪`: [u8(0xE8), 0x6D] // U+946A <cjk>
	`鈩`: [u8(0xE8), 0x6E] // U+9229 <cjk>
	`鑰`: [u8(0xE8), 0x6F] // U+9470 <cjk>
	`鑵`: [u8(0xE8), 0x70] // U+9475 <cjk>
	`鑷`: [u8(0xE8), 0x71] // U+9477 <cjk>
	`鑽`: [u8(0xE8), 0x72] // U+947D <cjk>
	`鑚`: [u8(0xE8), 0x73] // U+945A <cjk>
	`鑼`: [u8(0xE8), 0x74] // U+947C <cjk>
	`鑾`: [u8(0xE8), 0x75] // U+947E <cjk>
	`钁`: [u8(0xE8), 0x76] // U+9481 <cjk>
	`鑿`: [u8(0xE8), 0x77] // U+947F <cjk>
	`閂`: [u8(0xE8), 0x78] // U+9582 <cjk>
	`閇`: [u8(0xE8), 0x79] // U+9587 <cjk>
	`閊`: [u8(0xE8), 0x7A] // U+958A <cjk>
	`閔`: [u8(0xE8), 0x7B] // U+9594 <cjk>
	`閖`: [u8(0xE8), 0x7C] // U+9596 <cjk>
	`閘`: [u8(0xE8), 0x7D] // U+9598 <cjk>
	`閙`: [u8(0xE8), 0x7E] // U+9599 <cjk>
	`閠`: [u8(0xE8), 0x80] // U+95A0 <cjk>
	`閨`: [u8(0xE8), 0x81] // U+95A8 <cjk>
	`閧`: [u8(0xE8), 0x82] // U+95A7 <cjk>
	`閭`: [u8(0xE8), 0x83] // U+95AD <cjk>
	`閼`: [u8(0xE8), 0x84] // U+95BC <cjk>
	`閻`: [u8(0xE8), 0x85] // U+95BB <cjk>
	`閹`: [u8(0xE8), 0x86] // U+95B9 <cjk>
	`閾`: [u8(0xE8), 0x87] // U+95BE <cjk>
	`闊`: [u8(0xE8), 0x88] // U+95CA <cjk>
	`濶`: [u8(0xE8), 0x89] // U+6FF6 <cjk>
	`闃`: [u8(0xE8), 0x8A] // U+95C3 <cjk>
	`闍`: [u8(0xE8), 0x8B] // U+95CD <cjk>
	`闌`: [u8(0xE8), 0x8C] // U+95CC <cjk>
	`闕`: [u8(0xE8), 0x8D] // U+95D5 <cjk>
	`闔`: [u8(0xE8), 0x8E] // U+95D4 <cjk>
	`闖`: [u8(0xE8), 0x8F] // U+95D6 <cjk>
	`關`: [u8(0xE8), 0x90] // U+95DC <cjk>
	`闡`: [u8(0xE8), 0x91] // U+95E1 <cjk>
	`闥`: [u8(0xE8), 0x92] // U+95E5 <cjk>
	`闢`: [u8(0xE8), 0x93] // U+95E2 <cjk>
	`阡`: [u8(0xE8), 0x94] // U+9621 <cjk>
	`阨`: [u8(0xE8), 0x95] // U+9628 <cjk>
	`阮`: [u8(0xE8), 0x96] // U+962E <cjk>
	`阯`: [u8(0xE8), 0x97] // U+962F <cjk>
	`陂`: [u8(0xE8), 0x98] // U+9642 <cjk>
	`陌`: [u8(0xE8), 0x99] // U+964C <cjk>
	`陏`: [u8(0xE8), 0x9A] // U+964F <cjk>
	`陋`: [u8(0xE8), 0x9B] // U+964B <cjk>
	`陷`: [u8(0xE8), 0x9C] // U+9677 <cjk>
	`陜`: [u8(0xE8), 0x9D] // U+965C <cjk>
	`陞`: [u8(0xE8), 0x9E] // U+965E <cjk>
	`陝`: [u8(0xE8), 0x9F] // U+965D <cjk>
	`陟`: [u8(0xE8), 0xA0] // U+965F <cjk>
	`陦`: [u8(0xE8), 0xA1] // U+9666 <cjk>
	`陲`: [u8(0xE8), 0xA2] // U+9672 <cjk>
	`陬`: [u8(0xE8), 0xA3] // U+966C <cjk>
	`隍`: [u8(0xE8), 0xA4] // U+968D <cjk>
	`隘`: [u8(0xE8), 0xA5] // U+9698 <cjk>
	`隕`: [u8(0xE8), 0xA6] // U+9695 <cjk>
	`隗`: [u8(0xE8), 0xA7] // U+9697 <cjk>
	`險`: [u8(0xE8), 0xA8] // U+96AA <cjk>
	`隧`: [u8(0xE8), 0xA9] // U+96A7 <cjk>
	`隱`: [u8(0xE8), 0xAA] // U+96B1 <cjk>
	`隲`: [u8(0xE8), 0xAB] // U+96B2 <cjk>
	`隰`: [u8(0xE8), 0xAC] // U+96B0 <cjk>
	`隴`: [u8(0xE8), 0xAD] // U+96B4 <cjk>
	`隶`: [u8(0xE8), 0xAE] // U+96B6 <cjk>
	`隸`: [u8(0xE8), 0xAF] // U+96B8 <cjk>
	`隹`: [u8(0xE8), 0xB0] // U+96B9 <cjk>
	`雎`: [u8(0xE8), 0xB1] // U+96CE <cjk>
	`雋`: [u8(0xE8), 0xB2] // U+96CB <cjk>
	`雉`: [u8(0xE8), 0xB3] // U+96C9 <cjk>
	`雍`: [u8(0xE8), 0xB4] // U+96CD <cjk>
	`襍`: [u8(0xE8), 0xB5] // U+894D <cjk>
	`雜`: [u8(0xE8), 0xB6] // U+96DC <cjk>
	`霍`: [u8(0xE8), 0xB7] // U+970D <cjk>
	`雕`: [u8(0xE8), 0xB8] // U+96D5 <cjk>
	`雹`: [u8(0xE8), 0xB9] // U+96F9 <cjk>
	`霄`: [u8(0xE8), 0xBA] // U+9704 <cjk>
	`霆`: [u8(0xE8), 0xBB] // U+9706 <cjk>
	`霈`: [u8(0xE8), 0xBC] // U+9708 <cjk>
	`霓`: [u8(0xE8), 0xBD] // U+9713 <cjk>
	`霎`: [u8(0xE8), 0xBE] // U+970E <cjk>
	`霑`: [u8(0xE8), 0xBF] // U+9711 <cjk>
	`霏`: [u8(0xE8), 0xC0] // U+970F <cjk>
	`霖`: [u8(0xE8), 0xC1] // U+9716 <cjk>
	`霙`: [u8(0xE8), 0xC2] // U+9719 <cjk>
	`霤`: [u8(0xE8), 0xC3] // U+9724 <cjk>
	`霪`: [u8(0xE8), 0xC4] // U+972A <cjk>
	`霰`: [u8(0xE8), 0xC5] // U+9730 <cjk>
	`霹`: [u8(0xE8), 0xC6] // U+9739 <cjk>
	`霽`: [u8(0xE8), 0xC7] // U+973D <cjk>
	`霾`: [u8(0xE8), 0xC8] // U+973E <cjk>
	`靄`: [u8(0xE8), 0xC9] // U+9744 <cjk>
	`靆`: [u8(0xE8), 0xCA] // U+9746 <cjk>
	`靈`: [u8(0xE8), 0xCB] // U+9748 <cjk>
	`靂`: [u8(0xE8), 0xCC] // U+9742 <cjk>
	`靉`: [u8(0xE8), 0xCD] // U+9749 <cjk>
	`靜`: [u8(0xE8), 0xCE] // U+975C <cjk>
	`靠`: [u8(0xE8), 0xCF] // U+9760 <cjk>
	`靤`: [u8(0xE8), 0xD0] // U+9764 <cjk>
	`靦`: [u8(0xE8), 0xD1] // U+9766 <cjk>
	`靨`: [u8(0xE8), 0xD2] // U+9768 <cjk>
	`勒`: [u8(0xE8), 0xD3] // U+52D2 <cjk>
	`靫`: [u8(0xE8), 0xD4] // U+976B <cjk>
	`靱`: [u8(0xE8), 0xD5] // U+9771 <cjk>
	`靹`: [u8(0xE8), 0xD6] // U+9779 <cjk>
	`鞅`: [u8(0xE8), 0xD7] // U+9785 <cjk>
	`靼`: [u8(0xE8), 0xD8] // U+977C <cjk>
	`鞁`: [u8(0xE8), 0xD9] // U+9781 <cjk>
	`靺`: [u8(0xE8), 0xDA] // U+977A <cjk>
	`鞆`: [u8(0xE8), 0xDB] // U+9786 <cjk>
	`鞋`: [u8(0xE8), 0xDC] // U+978B <cjk>
	`鞏`: [u8(0xE8), 0xDD] // U+978F <cjk>
	`鞐`: [u8(0xE8), 0xDE] // U+9790 <cjk>
	`鞜`: [u8(0xE8), 0xDF] // U+979C <cjk>
	`鞨`: [u8(0xE8), 0xE0] // U+97A8 <cjk>
	`鞦`: [u8(0xE8), 0xE1] // U+97A6 <cjk>
	`鞣`: [u8(0xE8), 0xE2] // U+97A3 <cjk>
	`鞳`: [u8(0xE8), 0xE3] // U+97B3 <cjk>
	`鞴`: [u8(0xE8), 0xE4] // U+97B4 <cjk>
	`韃`: [u8(0xE8), 0xE5] // U+97C3 <cjk>
	`韆`: [u8(0xE8), 0xE6] // U+97C6 <cjk>
	`韈`: [u8(0xE8), 0xE7] // U+97C8 <cjk>
	`韋`: [u8(0xE8), 0xE8] // U+97CB <cjk>
	`韜`: [u8(0xE8), 0xE9] // U+97DC <cjk>
	`韭`: [u8(0xE8), 0xEA] // U+97ED <cjk>
	`齏`: [u8(0xE8), 0xEB] // U+9F4F <cjk>
	`韲`: [u8(0xE8), 0xEC] // U+97F2 <cjk>
	`竟`: [u8(0xE8), 0xED] // U+7ADF <cjk>
	`韶`: [u8(0xE8), 0xEE] // U+97F6 <cjk>
	`韵`: [u8(0xE8), 0xEF] // U+97F5 <cjk>
	`頏`: [u8(0xE8), 0xF0] // U+980F <cjk>
	`頌`: [u8(0xE8), 0xF1] // U+980C <cjk>
	`頸`: [u8(0xE8), 0xF2] // U+9838 <cjk>
	`頤`: [u8(0xE8), 0xF3] // U+9824 <cjk>
	`頡`: [u8(0xE8), 0xF4] // U+9821 <cjk>
	`頷`: [u8(0xE8), 0xF5] // U+9837 <cjk>
	`頽`: [u8(0xE8), 0xF6] // U+983D <cjk>
	`顆`: [u8(0xE8), 0xF7] // U+9846 <cjk>
	`顏`: [u8(0xE8), 0xF8] // U+984F <cjk>
	`顋`: [u8(0xE8), 0xF9] // U+984B <cjk>
	`顫`: [u8(0xE8), 0xFA] // U+986B <cjk>
	`顯`: [u8(0xE8), 0xFB] // U+986F <cjk>
	`顰`: [u8(0xE8), 0xFC] // U+9870 <cjk>
	`顱`: [u8(0xE9), 0x40] // U+9871 <cjk>
	`顴`: [u8(0xE9), 0x41] // U+9874 <cjk>
	`顳`: [u8(0xE9), 0x42] // U+9873 <cjk>
	`颪`: [u8(0xE9), 0x43] // U+98AA <cjk>
	`颯`: [u8(0xE9), 0x44] // U+98AF <cjk>
	`颱`: [u8(0xE9), 0x45] // U+98B1 <cjk>
	`颶`: [u8(0xE9), 0x46] // U+98B6 <cjk>
	`飄`: [u8(0xE9), 0x47] // U+98C4 <cjk>
	`飃`: [u8(0xE9), 0x48] // U+98C3 <cjk>
	`飆`: [u8(0xE9), 0x49] // U+98C6 <cjk>
	`飩`: [u8(0xE9), 0x4A] // U+98E9 <cjk>
	`飫`: [u8(0xE9), 0x4B] // U+98EB <cjk>
	`餃`: [u8(0xE9), 0x4C] // U+9903 <cjk>
	`餉`: [u8(0xE9), 0x4D] // U+9909 <cjk>
	`餒`: [u8(0xE9), 0x4E] // U+9912 <cjk>
	`餔`: [u8(0xE9), 0x4F] // U+9914 <cjk>
	`餘`: [u8(0xE9), 0x50] // U+9918 <cjk>
	`餡`: [u8(0xE9), 0x51] // U+9921 <cjk>
	`餝`: [u8(0xE9), 0x52] // U+991D <cjk>
	`餞`: [u8(0xE9), 0x53] // U+991E <cjk>
	`餤`: [u8(0xE9), 0x54] // U+9924 <cjk>
	`餠`: [u8(0xE9), 0x55] // U+9920 <cjk>
	`餬`: [u8(0xE9), 0x56] // U+992C <cjk>
	`餮`: [u8(0xE9), 0x57] // U+992E <cjk>
	`餽`: [u8(0xE9), 0x58] // U+993D <cjk>
	`餾`: [u8(0xE9), 0x59] // U+993E <cjk>
	`饂`: [u8(0xE9), 0x5A] // U+9942 <cjk>
	`饉`: [u8(0xE9), 0x5B] // U+9949 <cjk>
	`饅`: [u8(0xE9), 0x5C] // U+9945 <cjk>
	`饐`: [u8(0xE9), 0x5D] // U+9950 <cjk>
	`饋`: [u8(0xE9), 0x5E] // U+994B <cjk>
	`饑`: [u8(0xE9), 0x5F] // U+9951 <cjk>
	`饒`: [u8(0xE9), 0x60] // U+9952 <cjk>
	`饌`: [u8(0xE9), 0x61] // U+994C <cjk>
	`饕`: [u8(0xE9), 0x62] // U+9955 <cjk>
	`馗`: [u8(0xE9), 0x63] // U+9997 <cjk>
	`馘`: [u8(0xE9), 0x64] // U+9998 <cjk>
	`馥`: [u8(0xE9), 0x65] // U+99A5 <cjk>
	`馭`: [u8(0xE9), 0x66] // U+99AD <cjk>
	`馮`: [u8(0xE9), 0x67] // U+99AE <cjk>
	`馼`: [u8(0xE9), 0x68] // U+99BC <cjk>
	`駟`: [u8(0xE9), 0x69] // U+99DF <cjk>
	`駛`: [u8(0xE9), 0x6A] // U+99DB <cjk>
	`駝`: [u8(0xE9), 0x6B] // U+99DD <cjk>
	`駘`: [u8(0xE9), 0x6C] // U+99D8 <cjk>
	`駑`: [u8(0xE9), 0x6D] // U+99D1 <cjk>
	`駭`: [u8(0xE9), 0x6E] // U+99ED <cjk>
	`駮`: [u8(0xE9), 0x6F] // U+99EE <cjk>
	`駱`: [u8(0xE9), 0x70] // U+99F1 <cjk>
	`駲`: [u8(0xE9), 0x71] // U+99F2 <cjk>
	`駻`: [u8(0xE9), 0x72] // U+99FB <cjk>
	`駸`: [u8(0xE9), 0x73] // U+99F8 <cjk>
	`騁`: [u8(0xE9), 0x74] // U+9A01 <cjk>
	`騏`: [u8(0xE9), 0x75] // U+9A0F <cjk>
	`騅`: [u8(0xE9), 0x76] // U+9A05 <cjk>
	`駢`: [u8(0xE9), 0x77] // U+99E2 <cjk>
	`騙`: [u8(0xE9), 0x78] // U+9A19 <cjk>
	`騫`: [u8(0xE9), 0x79] // U+9A2B <cjk>
	`騷`: [u8(0xE9), 0x7A] // U+9A37 <cjk>
	`驅`: [u8(0xE9), 0x7B] // U+9A45 <cjk>
	`驂`: [u8(0xE9), 0x7C] // U+9A42 <cjk>
	`驀`: [u8(0xE9), 0x7D] // U+9A40 <cjk>
	`驃`: [u8(0xE9), 0x7E] // U+9A43 <cjk>
	`騾`: [u8(0xE9), 0x80] // U+9A3E <cjk>
	`驕`: [u8(0xE9), 0x81] // U+9A55 <cjk>
	`驍`: [u8(0xE9), 0x82] // U+9A4D <cjk>
	`驛`: [u8(0xE9), 0x83] // U+9A5B <cjk>
	`驗`: [u8(0xE9), 0x84] // U+9A57 <cjk>
	`驟`: [u8(0xE9), 0x85] // U+9A5F <cjk>
	`驢`: [u8(0xE9), 0x86] // U+9A62 <cjk>
	`驥`: [u8(0xE9), 0x87] // U+9A65 <cjk>
	`驤`: [u8(0xE9), 0x88] // U+9A64 <cjk>
	`驩`: [u8(0xE9), 0x89] // U+9A69 <cjk>
	`驫`: [u8(0xE9), 0x8A] // U+9A6B <cjk>
	`驪`: [u8(0xE9), 0x8B] // U+9A6A <cjk>
	`骭`: [u8(0xE9), 0x8C] // U+9AAD <cjk>
	`骰`: [u8(0xE9), 0x8D] // U+9AB0 <cjk>
	`骼`: [u8(0xE9), 0x8E] // U+9ABC <cjk>
	`髀`: [u8(0xE9), 0x8F] // U+9AC0 <cjk>
	`髏`: [u8(0xE9), 0x90] // U+9ACF <cjk>
	`髑`: [u8(0xE9), 0x91] // U+9AD1 <cjk>
	`髓`: [u8(0xE9), 0x92] // U+9AD3 <cjk>
	`體`: [u8(0xE9), 0x93] // U+9AD4 <cjk>
	`髞`: [u8(0xE9), 0x94] // U+9ADE <cjk>
	`髟`: [u8(0xE9), 0x95] // U+9ADF <cjk>
	`髢`: [u8(0xE9), 0x96] // U+9AE2 <cjk>
	`髣`: [u8(0xE9), 0x97] // U+9AE3 <cjk>
	`髦`: [u8(0xE9), 0x98] // U+9AE6 <cjk>
	`髯`: [u8(0xE9), 0x99] // U+9AEF <cjk>
	`髫`: [u8(0xE9), 0x9A] // U+9AEB <cjk>
	`髮`: [u8(0xE9), 0x9B] // U+9AEE <cjk>
	`髴`: [u8(0xE9), 0x9C] // U+9AF4 <cjk>
	`髱`: [u8(0xE9), 0x9D] // U+9AF1 <cjk>
	`髷`: [u8(0xE9), 0x9E] // U+9AF7 <cjk>
	`髻`: [u8(0xE9), 0x9F] // U+9AFB <cjk>
	`鬆`: [u8(0xE9), 0xA0] // U+9B06 <cjk>
	`鬘`: [u8(0xE9), 0xA1] // U+9B18 <cjk>
	`鬚`: [u8(0xE9), 0xA2] // U+9B1A <cjk>
	`鬟`: [u8(0xE9), 0xA3] // U+9B1F <cjk>
	`鬢`: [u8(0xE9), 0xA4] // U+9B22 <cjk>
	`鬣`: [u8(0xE9), 0xA5] // U+9B23 <cjk>
	`鬥`: [u8(0xE9), 0xA6] // U+9B25 <cjk>
	`鬧`: [u8(0xE9), 0xA7] // U+9B27 <cjk>
	`鬨`: [u8(0xE9), 0xA8] // U+9B28 <cjk>
	`鬩`: [u8(0xE9), 0xA9] // U+9B29 <cjk>
	`鬪`: [u8(0xE9), 0xAA] // U+9B2A <cjk>
	`鬮`: [u8(0xE9), 0xAB] // U+9B2E <cjk>
	`鬯`: [u8(0xE9), 0xAC] // U+9B2F <cjk>
	`鬲`: [u8(0xE9), 0xAD] // U+9B32 <cjk>
	`魄`: [u8(0xE9), 0xAE] // U+9B44 <cjk>
	`魃`: [u8(0xE9), 0xAF] // U+9B43 <cjk>
	`魏`: [u8(0xE9), 0xB0] // U+9B4F <cjk>
	`魍`: [u8(0xE9), 0xB1] // U+9B4D <cjk>
	`魎`: [u8(0xE9), 0xB2] // U+9B4E <cjk>
	`魑`: [u8(0xE9), 0xB3] // U+9B51 <cjk>
	`魘`: [u8(0xE9), 0xB4] // U+9B58 <cjk>
	`魴`: [u8(0xE9), 0xB5] // U+9B74 <cjk>
	`鮓`: [u8(0xE9), 0xB6] // U+9B93 <cjk>
	`鮃`: [u8(0xE9), 0xB7] // U+9B83 <cjk>
	`鮑`: [u8(0xE9), 0xB8] // U+9B91 <cjk>
	`鮖`: [u8(0xE9), 0xB9] // U+9B96 <cjk>
	`鮗`: [u8(0xE9), 0xBA] // U+9B97 <cjk>
	`鮟`: [u8(0xE9), 0xBB] // U+9B9F <cjk>
	`鮠`: [u8(0xE9), 0xBC] // U+9BA0 <cjk>
	`鮨`: [u8(0xE9), 0xBD] // U+9BA8 <cjk>
	`鮴`: [u8(0xE9), 0xBE] // U+9BB4 <cjk>
	`鯀`: [u8(0xE9), 0xBF] // U+9BC0 <cjk>
	`鯊`: [u8(0xE9), 0xC0] // U+9BCA <cjk>
	`鮹`: [u8(0xE9), 0xC1] // U+9BB9 <cjk>
	`鯆`: [u8(0xE9), 0xC2] // U+9BC6 <cjk>
	`鯏`: [u8(0xE9), 0xC3] // U+9BCF <cjk>
	`鯑`: [u8(0xE9), 0xC4] // U+9BD1 <cjk>
	`鯒`: [u8(0xE9), 0xC5] // U+9BD2 <cjk>
	`鯣`: [u8(0xE9), 0xC6] // U+9BE3 <cjk>
	`鯢`: [u8(0xE9), 0xC7] // U+9BE2 <cjk>
	`鯤`: [u8(0xE9), 0xC8] // U+9BE4 <cjk>
	`鯔`: [u8(0xE9), 0xC9] // U+9BD4 <cjk>
	`鯡`: [u8(0xE9), 0xCA] // U+9BE1 <cjk>
	`鰺`: [u8(0xE9), 0xCB] // U+9C3A <cjk>
	`鯲`: [u8(0xE9), 0xCC] // U+9BF2 <cjk>
	`鯱`: [u8(0xE9), 0xCD] // U+9BF1 <cjk>
	`鯰`: [u8(0xE9), 0xCE] // U+9BF0 <cjk>
	`鰕`: [u8(0xE9), 0xCF] // U+9C15 <cjk>
	`鰔`: [u8(0xE9), 0xD0] // U+9C14 <cjk>
	`鰉`: [u8(0xE9), 0xD1] // U+9C09 <cjk>
	`鰓`: [u8(0xE9), 0xD2] // U+9C13 <cjk>
	`鰌`: [u8(0xE9), 0xD3] // U+9C0C <cjk>
	`鰆`: [u8(0xE9), 0xD4] // U+9C06 <cjk>
	`鰈`: [u8(0xE9), 0xD5] // U+9C08 <cjk>
	`鰒`: [u8(0xE9), 0xD6] // U+9C12 <cjk>
	`鰊`: [u8(0xE9), 0xD7] // U+9C0A <cjk>
	`鰄`: [u8(0xE9), 0xD8] // U+9C04 <cjk>
	`鰮`: [u8(0xE9), 0xD9] // U+9C2E <cjk>
	`鰛`: [u8(0xE9), 0xDA] // U+9C1B <cjk>
	`鰥`: [u8(0xE9), 0xDB] // U+9C25 <cjk>
	`鰤`: [u8(0xE9), 0xDC] // U+9C24 <cjk>
	`鰡`: [u8(0xE9), 0xDD] // U+9C21 <cjk>
	`鰰`: [u8(0xE9), 0xDE] // U+9C30 <cjk>
	`鱇`: [u8(0xE9), 0xDF] // U+9C47 <cjk>
	`鰲`: [u8(0xE9), 0xE0] // U+9C32 <cjk>
	`鱆`: [u8(0xE9), 0xE1] // U+9C46 <cjk>
	`鰾`: [u8(0xE9), 0xE2] // U+9C3E <cjk>
	`鱚`: [u8(0xE9), 0xE3] // U+9C5A <cjk>
	`鱠`: [u8(0xE9), 0xE4] // U+9C60 <cjk>
	`鱧`: [u8(0xE9), 0xE5] // U+9C67 <cjk>
	`鱶`: [u8(0xE9), 0xE6] // U+9C76 <cjk>
	`鱸`: [u8(0xE9), 0xE7] // U+9C78 <cjk>
	`鳧`: [u8(0xE9), 0xE8] // U+9CE7 <cjk>
	`鳬`: [u8(0xE9), 0xE9] // U+9CEC <cjk>
	`鳰`: [u8(0xE9), 0xEA] // U+9CF0 <cjk>
	`鴉`: [u8(0xE9), 0xEB] // U+9D09 <cjk>
	`鴈`: [u8(0xE9), 0xEC] // U+9D08 <cjk>
	`鳫`: [u8(0xE9), 0xED] // U+9CEB <cjk>
	`鴃`: [u8(0xE9), 0xEE] // U+9D03 <cjk>
	`鴆`: [u8(0xE9), 0xEF] // U+9D06 <cjk>
	`鴪`: [u8(0xE9), 0xF0] // U+9D2A <cjk>
	`鴦`: [u8(0xE9), 0xF1] // U+9D26 <cjk>
	`鶯`: [u8(0xE9), 0xF2] // U+9DAF <cjk>
	`鴣`: [u8(0xE9), 0xF3] // U+9D23 <cjk>
	`鴟`: [u8(0xE9), 0xF4] // U+9D1F <cjk>
	`鵄`: [u8(0xE9), 0xF5] // U+9D44 <cjk>
	`鴕`: [u8(0xE9), 0xF6] // U+9D15 <cjk>
	`鴒`: [u8(0xE9), 0xF7] // U+9D12 <cjk>
	`鵁`: [u8(0xE9), 0xF8] // U+9D41 <cjk>
	`鴿`: [u8(0xE9), 0xF9] // U+9D3F <cjk>
	`鴾`: [u8(0xE9), 0xFA] // U+9D3E <cjk>
	`鵆`: [u8(0xE9), 0xFB] // U+9D46 <cjk>
	`鵈`: [u8(0xE9), 0xFC] // U+9D48 <cjk>
	`鵝`: [u8(0xEA), 0x40] // U+9D5D <cjk>
	`鵞`: [u8(0xEA), 0x41] // U+9D5E <cjk>
	`鵤`: [u8(0xEA), 0x42] // U+9D64 <cjk>
	`鵑`: [u8(0xEA), 0x43] // U+9D51 <cjk>
	`鵐`: [u8(0xEA), 0x44] // U+9D50 <cjk>
	`鵙`: [u8(0xEA), 0x45] // U+9D59 <cjk>
	`鵲`: [u8(0xEA), 0x46] // U+9D72 <cjk>
	`鶉`: [u8(0xEA), 0x47] // U+9D89 <cjk>
	`鶇`: [u8(0xEA), 0x48] // U+9D87 <cjk>
	`鶫`: [u8(0xEA), 0x49] // U+9DAB <cjk>
	`鵯`: [u8(0xEA), 0x4A] // U+9D6F <cjk>
	`鵺`: [u8(0xEA), 0x4B] // U+9D7A <cjk>
	`鶚`: [u8(0xEA), 0x4C] // U+9D9A <cjk>
	`鶤`: [u8(0xEA), 0x4D] // U+9DA4 <cjk>
	`鶩`: [u8(0xEA), 0x4E] // U+9DA9 <cjk>
	`鶲`: [u8(0xEA), 0x4F] // U+9DB2 <cjk>
	`鷄`: [u8(0xEA), 0x50] // U+9DC4 <cjk>
	`鷁`: [u8(0xEA), 0x51] // U+9DC1 <cjk>
	`鶻`: [u8(0xEA), 0x52] // U+9DBB <cjk>
	`鶸`: [u8(0xEA), 0x53] // U+9DB8 <cjk>
	`鶺`: [u8(0xEA), 0x54] // U+9DBA <cjk>
	`鷆`: [u8(0xEA), 0x55] // U+9DC6 <cjk>
	`鷏`: [u8(0xEA), 0x56] // U+9DCF <cjk>
	`鷂`: [u8(0xEA), 0x57] // U+9DC2 <cjk>
	`鷙`: [u8(0xEA), 0x58] // U+9DD9 <cjk>
	`鷓`: [u8(0xEA), 0x59] // U+9DD3 <cjk>
	`鷸`: [u8(0xEA), 0x5A] // U+9DF8 <cjk>
	`鷦`: [u8(0xEA), 0x5B] // U+9DE6 <cjk>
	`鷭`: [u8(0xEA), 0x5C] // U+9DED <cjk>
	`鷯`: [u8(0xEA), 0x5D] // U+9DEF <cjk>
	`鷽`: [u8(0xEA), 0x5E] // U+9DFD <cjk>
	`鸚`: [u8(0xEA), 0x5F] // U+9E1A <cjk>
	`鸛`: [u8(0xEA), 0x60] // U+9E1B <cjk>
	`鸞`: [u8(0xEA), 0x61] // U+9E1E <cjk>
	`鹵`: [u8(0xEA), 0x62] // U+9E75 <cjk>
	`鹹`: [u8(0xEA), 0x63] // U+9E79 <cjk>
	`鹽`: [u8(0xEA), 0x64] // U+9E7D <cjk>
	`麁`: [u8(0xEA), 0x65] // U+9E81 <cjk>
	`麈`: [u8(0xEA), 0x66] // U+9E88 <cjk>
	`麋`: [u8(0xEA), 0x67] // U+9E8B <cjk>
	`麌`: [u8(0xEA), 0x68] // U+9E8C <cjk>
	`麒`: [u8(0xEA), 0x69] // U+9E92 <cjk>
	`麕`: [u8(0xEA), 0x6A] // U+9E95 <cjk>
	`麑`: [u8(0xEA), 0x6B] // U+9E91 <cjk>
	`麝`: [u8(0xEA), 0x6C] // U+9E9D <cjk>
	`麥`: [u8(0xEA), 0x6D] // U+9EA5 <cjk>
	`麩`: [u8(0xEA), 0x6E] // U+9EA9 <cjk>
	`麸`: [u8(0xEA), 0x6F] // U+9EB8 <cjk>
	`麪`: [u8(0xEA), 0x70] // U+9EAA <cjk>
	`麭`: [u8(0xEA), 0x71] // U+9EAD <cjk>
	`靡`: [u8(0xEA), 0x72] // U+9761 <cjk>
	`黌`: [u8(0xEA), 0x73] // U+9ECC <cjk>
	`黎`: [u8(0xEA), 0x74] // U+9ECE <cjk>
	`黏`: [u8(0xEA), 0x75] // U+9ECF <cjk>
	`黐`: [u8(0xEA), 0x76] // U+9ED0 <cjk>
	`黔`: [u8(0xEA), 0x77] // U+9ED4 <cjk>
	`黜`: [u8(0xEA), 0x78] // U+9EDC <cjk>
	`點`: [u8(0xEA), 0x79] // U+9EDE <cjk>
	`黝`: [u8(0xEA), 0x7A] // U+9EDD <cjk>
	`黠`: [u8(0xEA), 0x7B] // U+9EE0 <cjk>
	`黥`: [u8(0xEA), 0x7C] // U+9EE5 <cjk>
	`黨`: [u8(0xEA), 0x7D] // U+9EE8 <cjk>
	`黯`: [u8(0xEA), 0x7E] // U+9EEF <cjk>
	`黴`: [u8(0xEA), 0x80] // U+9EF4 <cjk>
	`黶`: [u8(0xEA), 0x81] // U+9EF6 <cjk>
	`黷`: [u8(0xEA), 0x82] // U+9EF7 <cjk>
	`黹`: [u8(0xEA), 0x83] // U+9EF9 <cjk>
	`黻`: [u8(0xEA), 0x84] // U+9EFB <cjk>
	`黼`: [u8(0xEA), 0x85] // U+9EFC <cjk>
	`黽`: [u8(0xEA), 0x86] // U+9EFD <cjk>
	`鼇`: [u8(0xEA), 0x87] // U+9F07 <cjk>
	`鼈`: [u8(0xEA), 0x88] // U+9F08 <cjk>
	`皷`: [u8(0xEA), 0x89] // U+76B7 <cjk>
	`鼕`: [u8(0xEA), 0x8A] // U+9F15 <cjk>
	`鼡`: [u8(0xEA), 0x8B] // U+9F21 <cjk>
	`鼬`: [u8(0xEA), 0x8C] // U+9F2C <cjk>
	`鼾`: [u8(0xEA), 0x8D] // U+9F3E <cjk>
	`齊`: [u8(0xEA), 0x8E] // U+9F4A <cjk>
	`齒`: [u8(0xEA), 0x8F] // U+9F52 <cjk>
	`齔`: [u8(0xEA), 0x90] // U+9F54 <cjk>
	`齣`: [u8(0xEA), 0x91] // U+9F63 <cjk>
	`齟`: [u8(0xEA), 0x92] // U+9F5F <cjk>
	`齠`: [u8(0xEA), 0x93] // U+9F60 <cjk>
	`齡`: [u8(0xEA), 0x94] // U+9F61 <cjk>
	`齦`: [u8(0xEA), 0x95] // U+9F66 <cjk>
	`齧`: [u8(0xEA), 0x96] // U+9F67 <cjk>
	`齬`: [u8(0xEA), 0x97] // U+9F6C <cjk>
	`齪`: [u8(0xEA), 0x98] // U+9F6A <cjk>
	`齷`: [u8(0xEA), 0x99] // U+9F77 <cjk>
	`齲`: [u8(0xEA), 0x9A] // U+9F72 <cjk>
	`齶`: [u8(0xEA), 0x9B] // U+9F76 <cjk>
	`龕`: [u8(0xEA), 0x9C] // U+9F95 <cjk>
	`龜`: [u8(0xEA), 0x9D] // U+9F9C <cjk>
	`龠`: [u8(0xEA), 0x9E] // U+9FA0 <cjk>
	`堯`: [u8(0xEA), 0x9F] // U+582F <cjk>
	`槇`: [u8(0xEA), 0xA0] // U+69C7 <cjk>
	`遙`: [u8(0xEA), 0xA1] // U+9059 <cjk>
	`瑤`: [u8(0xEA), 0xA2] // U+7464 <cjk>
	`凜`: [u8(0xEA), 0xA3] // U+51DC <cjk>
	`熙`: [u8(0xEA), 0xA4] // U+7199 <cjk>
	`噓`: [u8(0xEA), 0xA5] // U+5653 <cjk>
	`巢`: [u8(0xEA), 0xA6] // U+5DE2 <cjk>
	`帔`: [u8(0xEA), 0xA7] // U+5E14 <cjk>
	`帘`: [u8(0xEA), 0xA8] // U+5E18 <cjk>
	`幘`: [u8(0xEA), 0xA9] // U+5E58 <cjk>
	`幞`: [u8(0xEA), 0xAA] // U+5E5E <cjk>
	`庾`: [u8(0xEA), 0xAB] // U+5EBE <cjk>
	`廊`: [u8(0xEA), 0xAC] // U+F928 CJK COMPATIBILITY IDEOGRAPH-F928
	`廋`: [u8(0xEA), 0xAD] // U+5ECB <cjk>
	`廹`: [u8(0xEA), 0xAE] // U+5EF9 <cjk>
	`开`: [u8(0xEA), 0xAF] // U+5F00 <cjk>
	`异`: [u8(0xEA), 0xB0] // U+5F02 <cjk>
	`弇`: [u8(0xEA), 0xB1] // U+5F07 <cjk>
	`弝`: [u8(0xEA), 0xB2] // U+5F1D <cjk>
	`弣`: [u8(0xEA), 0xB3] // U+5F23 <cjk>
	`弴`: [u8(0xEA), 0xB4] // U+5F34 <cjk>
	`弶`: [u8(0xEA), 0xB5] // U+5F36 <cjk>
	`弽`: [u8(0xEA), 0xB6] // U+5F3D <cjk>
	`彀`: [u8(0xEA), 0xB7] // U+5F40 <cjk>
	`彅`: [u8(0xEA), 0xB8] // U+5F45 <cjk>
	`彔`: [u8(0xEA), 0xB9] // U+5F54 <cjk>
	`彘`: [u8(0xEA), 0xBA] // U+5F58 <cjk>
	`彤`: [u8(0xEA), 0xBB] // U+5F64 <cjk>
	`彧`: [u8(0xEA), 0xBC] // U+5F67 <cjk>
	`彽`: [u8(0xEA), 0xBD] // U+5F7D <cjk>
	`徉`: [u8(0xEA), 0xBE] // U+5F89 <cjk>
	`徜`: [u8(0xEA), 0xBF] // U+5F9C <cjk>
	`徧`: [u8(0xEA), 0xC0] // U+5FA7 <cjk>
	`徯`: [u8(0xEA), 0xC1] // U+5FAF <cjk>
	`徵`: [u8(0xEA), 0xC2] // U+5FB5 <cjk>
	`德`: [u8(0xEA), 0xC3] // U+5FB7 <cjk>
	`忉`: [u8(0xEA), 0xC4] // U+5FC9 <cjk>
	`忞`: [u8(0xEA), 0xC5] // U+5FDE <cjk>
	`忡`: [u8(0xEA), 0xC6] // U+5FE1 <cjk>
	`忩`: [u8(0xEA), 0xC7] // U+5FE9 <cjk>
	`怍`: [u8(0xEA), 0xC8] // U+600D <cjk>
	`怔`: [u8(0xEA), 0xC9] // U+6014 <cjk>
	`怘`: [u8(0xEA), 0xCA] // U+6018 <cjk>
	`怳`: [u8(0xEA), 0xCB] // U+6033 <cjk>
	`怵`: [u8(0xEA), 0xCC] // U+6035 <cjk>
	`恇`: [u8(0xEA), 0xCD] // U+6047 <cjk>
	`悔`: [u8(0xEA), 0xCE] // U+FA3D CJK COMPATIBILITY IDEOGRAPH-FA3D
	`悝`: [u8(0xEA), 0xCF] // U+609D <cjk>
	`悞`: [u8(0xEA), 0xD0] // U+609E <cjk>
	`惋`: [u8(0xEA), 0xD1] // U+60CB <cjk>
	`惔`: [u8(0xEA), 0xD2] // U+60D4 <cjk>
	`惕`: [u8(0xEA), 0xD3] // U+60D5 <cjk>
	`惝`: [u8(0xEA), 0xD4] // U+60DD <cjk>
	`惸`: [u8(0xEA), 0xD5] // U+60F8 <cjk>
	`愜`: [u8(0xEA), 0xD6] // U+611C <cjk>
	`愫`: [u8(0xEA), 0xD7] // U+612B <cjk>
	`愰`: [u8(0xEA), 0xD8] // U+6130 <cjk>
	`愷`: [u8(0xEA), 0xD9] // U+6137 <cjk>
	`慨`: [u8(0xEA), 0xDA] // U+FA3E CJK COMPATIBILITY IDEOGRAPH-FA3E
	`憍`: [u8(0xEA), 0xDB] // U+618D <cjk>
	`憎`: [u8(0xEA), 0xDC] // U+FA3F CJK COMPATIBILITY IDEOGRAPH-FA3F
	`憼`: [u8(0xEA), 0xDD] // U+61BC <cjk>
	`憹`: [u8(0xEA), 0xDE] // U+61B9 <cjk>
	`懲`: [u8(0xEA), 0xDF] // U+FA40 CJK COMPATIBILITY IDEOGRAPH-FA40
	`戢`: [u8(0xEA), 0xE0] // U+6222 <cjk>
	`戾`: [u8(0xEA), 0xE1] // U+623E <cjk>
	`扃`: [u8(0xEA), 0xE2] // U+6243 <cjk>
	`扖`: [u8(0xEA), 0xE3] // U+6256 <cjk>
	`扚`: [u8(0xEA), 0xE4] // U+625A <cjk>
	`扯`: [u8(0xEA), 0xE5] // U+626F <cjk>
	`抅`: [u8(0xEA), 0xE6] // U+6285 <cjk>
	`拄`: [u8(0xEA), 0xE7] // U+62C4 <cjk>
	`拖`: [u8(0xEA), 0xE8] // U+62D6 <cjk>
	`拼`: [u8(0xEA), 0xE9] // U+62FC <cjk>
	`挊`: [u8(0xEA), 0xEA] // U+630A <cjk>
	`挘`: [u8(0xEA), 0xEB] // U+6318 <cjk>
	`挹`: [u8(0xEA), 0xEC] // U+6339 <cjk>
	`捃`: [u8(0xEA), 0xED] // U+6343 <cjk>
	`捥`: [u8(0xEA), 0xEE] // U+6365 <cjk>
	`捼`: [u8(0xEA), 0xEF] // U+637C <cjk>
	`揥`: [u8(0xEA), 0xF0] // U+63E5 <cjk>
	`揭`: [u8(0xEA), 0xF1] // U+63ED <cjk>
	`揵`: [u8(0xEA), 0xF2] // U+63F5 <cjk>
	`搐`: [u8(0xEA), 0xF3] // U+6410 <cjk>
	`搔`: [u8(0xEA), 0xF4] // U+6414 <cjk>
	`搢`: [u8(0xEA), 0xF5] // U+6422 <cjk>
	`摹`: [u8(0xEA), 0xF6] // U+6479 <cjk>
	`摑`: [u8(0xEA), 0xF7] // U+6451 <cjk>
	`摠`: [u8(0xEA), 0xF8] // U+6460 <cjk>
	`摭`: [u8(0xEA), 0xF9] // U+646D <cjk>
	`擎`: [u8(0xEA), 0xFA] // U+64CE <cjk>
	`撾`: [u8(0xEA), 0xFB] // U+64BE <cjk>
	`撿`: [u8(0xEA), 0xFC] // U+64BF <cjk>
	`擄`: [u8(0xEB), 0x40] // U+64C4 <cjk>
	`擊`: [u8(0xEB), 0x41] // U+64CA <cjk>
	`擐`: [u8(0xEB), 0x42] // U+64D0 <cjk>
	`擷`: [u8(0xEB), 0x43] // U+64F7 <cjk>
	`擻`: [u8(0xEB), 0x44] // U+64FB <cjk>
	`攢`: [u8(0xEB), 0x45] // U+6522 <cjk>
	`攩`: [u8(0xEB), 0x46] // U+6529 <cjk>
	`敏`: [u8(0xEB), 0x47] // U+FA41 CJK COMPATIBILITY IDEOGRAPH-FA41
	`敧`: [u8(0xEB), 0x48] // U+6567 <cjk>
	`斝`: [u8(0xEB), 0x49] // U+659D <cjk>
	`既`: [u8(0xEB), 0x4A] // U+FA42 CJK COMPATIBILITY IDEOGRAPH-FA42
	`昀`: [u8(0xEB), 0x4B] // U+6600 <cjk>
	`昉`: [u8(0xEB), 0x4C] // U+6609 <cjk>
	`昕`: [u8(0xEB), 0x4D] // U+6615 <cjk>
	`昞`: [u8(0xEB), 0x4E] // U+661E <cjk>
	`昺`: [u8(0xEB), 0x4F] // U+663A <cjk>
	`昢`: [u8(0xEB), 0x50] // U+6622 <cjk>
	`昤`: [u8(0xEB), 0x51] // U+6624 <cjk>
	`昫`: [u8(0xEB), 0x52] // U+662B <cjk>
	`昰`: [u8(0xEB), 0x53] // U+6630 <cjk>
	`昱`: [u8(0xEB), 0x54] // U+6631 <cjk>
	`昳`: [u8(0xEB), 0x55] // U+6633 <cjk>
	`曻`: [u8(0xEB), 0x56] // U+66FB <cjk>
	`晈`: [u8(0xEB), 0x57] // U+6648 <cjk>
	`晌`: [u8(0xEB), 0x58] // U+664C <cjk>
	`𣇄`: [u8(0xEB), 0x59] // U+231C4 <cjk>
	`晙`: [u8(0xEB), 0x5A] // U+6659 <cjk>
	`晚`: [u8(0xEB), 0x5B] // U+665A <cjk>
	`晡`: [u8(0xEB), 0x5C] // U+6661 <cjk>
	`晥`: [u8(0xEB), 0x5D] // U+6665 <cjk>
	`晳`: [u8(0xEB), 0x5E] // U+6673 <cjk>
	`晷`: [u8(0xEB), 0x5F] // U+6677 <cjk>
	`晸`: [u8(0xEB), 0x60] // U+6678 <cjk>
	`暍`: [u8(0xEB), 0x61] // U+668D <cjk>
	`暑`: [u8(0xEB), 0x62] // U+FA43 CJK COMPATIBILITY IDEOGRAPH-FA43
	`暠`: [u8(0xEB), 0x63] // U+66A0 <cjk>
	`暲`: [u8(0xEB), 0x64] // U+66B2 <cjk>
	`暻`: [u8(0xEB), 0x65] // U+66BB <cjk>
	`曆`: [u8(0xEB), 0x66] // U+66C6 <cjk>
	`曈`: [u8(0xEB), 0x67] // U+66C8 <cjk>
	`㬢`: [u8(0xEB), 0x68] // U+3B22 <cjk>
	`曛`: [u8(0xEB), 0x69] // U+66DB <cjk>
	`曨`: [u8(0xEB), 0x6A] // U+66E8 <cjk>
	`曺`: [u8(0xEB), 0x6B] // U+66FA <cjk>
	`朓`: [u8(0xEB), 0x6C] // U+6713 <cjk>
	`朗`: [u8(0xEB), 0x6D] // U+F929 CJK COMPATIBILITY IDEOGRAPH-F929
	`朳`: [u8(0xEB), 0x6E] // U+6733 <cjk>
	`杦`: [u8(0xEB), 0x6F] // U+6766 <cjk>
	`杇`: [u8(0xEB), 0x70] // U+6747 <cjk>
	`杈`: [u8(0xEB), 0x71] // U+6748 <cjk>
	`杻`: [u8(0xEB), 0x72] // U+677B <cjk>
	`极`: [u8(0xEB), 0x73] // U+6781 <cjk>
	`枓`: [u8(0xEB), 0x74] // U+6793 <cjk>
	`枘`: [u8(0xEB), 0x75] // U+6798 <cjk>
	`枛`: [u8(0xEB), 0x76] // U+679B <cjk>
	`枻`: [u8(0xEB), 0x77] // U+67BB <cjk>
	`柹`: [u8(0xEB), 0x78] // U+67F9 <cjk>
	`柀`: [u8(0xEB), 0x79] // U+67C0 <cjk>
	`柗`: [u8(0xEB), 0x7A] // U+67D7 <cjk>
	`柼`: [u8(0xEB), 0x7B] // U+67FC <cjk>
	`栁`: [u8(0xEB), 0x7C] // U+6801 <cjk>
	`桒`: [u8(0xEB), 0x7D] // U+6852 <cjk>
	`栝`: [u8(0xEB), 0x7E] // U+681D <cjk>
	`栬`: [u8(0xEB), 0x80] // U+682C <cjk>
	`栱`: [u8(0xEB), 0x81] // U+6831 <cjk>
	`桛`: [u8(0xEB), 0x82] // U+685B <cjk>
	`桲`: [u8(0xEB), 0x83] // U+6872 <cjk>
	`桵`: [u8(0xEB), 0x84] // U+6875 <cjk>
	`梅`: [u8(0xEB), 0x85] // U+FA44 CJK COMPATIBILITY IDEOGRAPH-FA44
	`梣`: [u8(0xEB), 0x86] // U+68A3 <cjk>
	`梥`: [u8(0xEB), 0x87] // U+68A5 <cjk>
	`梲`: [u8(0xEB), 0x88] // U+68B2 <cjk>
	`棈`: [u8(0xEB), 0x89] // U+68C8 <cjk>
	`棐`: [u8(0xEB), 0x8A] // U+68D0 <cjk>
	`棨`: [u8(0xEB), 0x8B] // U+68E8 <cjk>
	`棭`: [u8(0xEB), 0x8C] // U+68ED <cjk>
	`棰`: [u8(0xEB), 0x8D] // U+68F0 <cjk>
	`棱`: [u8(0xEB), 0x8E] // U+68F1 <cjk>
	`棼`: [u8(0xEB), 0x8F] // U+68FC <cjk>
	`椊`: [u8(0xEB), 0x90] // U+690A <cjk>
	`楉`: [u8(0xEB), 0x91] // U+6949 <cjk>
	`𣗄`: [u8(0xEB), 0x92] // U+235C4 <cjk>
	`椵`: [u8(0xEB), 0x93] // U+6935 <cjk>
	`楂`: [u8(0xEB), 0x94] // U+6942 <cjk>
	`楗`: [u8(0xEB), 0x95] // U+6957 <cjk>
	`楣`: [u8(0xEB), 0x96] // U+6963 <cjk>
	`楤`: [u8(0xEB), 0x97] // U+6964 <cjk>
	`楨`: [u8(0xEB), 0x98] // U+6968 <cjk>
	`榀`: [u8(0xEB), 0x99] // U+6980 <cjk>
	`﨔`: [u8(0xEB), 0x9A] // U+FA14 CJK COMPATIBILITY IDEOGRAPH-FA14
	`榥`: [u8(0xEB), 0x9B] // U+69A5 <cjk>
	`榭`: [u8(0xEB), 0x9C] // U+69AD <cjk>
	`槏`: [u8(0xEB), 0x9D] // U+69CF <cjk>
	`㮶`: [u8(0xEB), 0x9E] // U+3BB6 <cjk>
	`㯃`: [u8(0xEB), 0x9F] // U+3BC3 <cjk>
	`槢`: [u8(0xEB), 0xA0] // U+69E2 <cjk>
	`槩`: [u8(0xEB), 0xA1] // U+69E9 <cjk>
	`槪`: [u8(0xEB), 0xA2] // U+69EA <cjk>
	`槵`: [u8(0xEB), 0xA3] // U+69F5 <cjk>
	`槶`: [u8(0xEB), 0xA4] // U+69F6 <cjk>
	`樏`: [u8(0xEB), 0xA5] // U+6A0F <cjk>
	`樕`: [u8(0xEB), 0xA6] // U+6A15 <cjk>
	`𣜿`: [u8(0xEB), 0xA7] // U+2373F <cjk>
	`樻`: [u8(0xEB), 0xA8] // U+6A3B <cjk>
	`樾`: [u8(0xEB), 0xA9] // U+6A3E <cjk>
	`橅`: [u8(0xEB), 0xAA] // U+6A45 <cjk>
	`橐`: [u8(0xEB), 0xAB] // U+6A50 <cjk>
	`橖`: [u8(0xEB), 0xAC] // U+6A56 <cjk>
	`橛`: [u8(0xEB), 0xAD] // U+6A5B <cjk>
	`橫`: [u8(0xEB), 0xAE] // U+6A6B <cjk>
	`橳`: [u8(0xEB), 0xAF] // U+6A73 <cjk>
	`𣝣`: [u8(0xEB), 0xB0] // U+23763 <cjk>
	`檉`: [u8(0xEB), 0xB1] // U+6A89 <cjk>
	`檔`: [u8(0xEB), 0xB2] // U+6A94 <cjk>
	`檝`: [u8(0xEB), 0xB3] // U+6A9D <cjk>
	`檞`: [u8(0xEB), 0xB4] // U+6A9E <cjk>
	`檥`: [u8(0xEB), 0xB5] // U+6AA5 <cjk>
	`櫤`: [u8(0xEB), 0xB6] // U+6AE4 <cjk>
	`櫧`: [u8(0xEB), 0xB7] // U+6AE7 <cjk>
	`㰏`: [u8(0xEB), 0xB8] // U+3C0F <cjk>
	`欄`: [u8(0xEB), 0xB9] // U+F91D CJK COMPATIBILITY IDEOGRAPH-F91D
	`欛`: [u8(0xEB), 0xBA] // U+6B1B <cjk>
	`欞`: [u8(0xEB), 0xBB] // U+6B1E <cjk>
	`欬`: [u8(0xEB), 0xBC] // U+6B2C <cjk>
	`欵`: [u8(0xEB), 0xBD] // U+6B35 <cjk>
	`歆`: [u8(0xEB), 0xBE] // U+6B46 <cjk>
	`歖`: [u8(0xEB), 0xBF] // U+6B56 <cjk>
	`歠`: [u8(0xEB), 0xC0] // U+6B60 <cjk>
	`步`: [u8(0xEB), 0xC1] // U+6B65 <cjk>
	`歧`: [u8(0xEB), 0xC2] // U+6B67 <cjk>
	`歷`: [u8(0xEB), 0xC3] // U+6B77 <cjk>
	`殂`: [u8(0xEB), 0xC4] // U+6B82 <cjk>
	`殩`: [u8(0xEB), 0xC5] // U+6BA9 <cjk>
	`殭`: [u8(0xEB), 0xC6] // U+6BAD <cjk>
	`殺`: [u8(0xEB), 0xC7] // U+F970 CJK COMPATIBILITY IDEOGRAPH-F970
	`每`: [u8(0xEB), 0xC8] // U+6BCF <cjk>
	`毖`: [u8(0xEB), 0xC9] // U+6BD6 <cjk>
	`毗`: [u8(0xEB), 0xCA] // U+6BD7 <cjk>
	`毿`: [u8(0xEB), 0xCB] // U+6BFF <cjk>
	`氅`: [u8(0xEB), 0xCC] // U+6C05 <cjk>
	`氐`: [u8(0xEB), 0xCD] // U+6C10 <cjk>
	`氳`: [u8(0xEB), 0xCE] // U+6C33 <cjk>
	`汙`: [u8(0xEB), 0xCF] // U+6C59 <cjk>
	`汜`: [u8(0xEB), 0xD0] // U+6C5C <cjk>
	`沪`: [u8(0xEB), 0xD1] // U+6CAA <cjk>
	`汴`: [u8(0xEB), 0xD2] // U+6C74 <cjk>
	`汶`: [u8(0xEB), 0xD3] // U+6C76 <cjk>
	`沅`: [u8(0xEB), 0xD4] // U+6C85 <cjk>
	`沆`: [u8(0xEB), 0xD5] // U+6C86 <cjk>
	`沘`: [u8(0xEB), 0xD6] // U+6C98 <cjk>
	`沜`: [u8(0xEB), 0xD7] // U+6C9C <cjk>
	`泻`: [u8(0xEB), 0xD8] // U+6CFB <cjk>
	`泆`: [u8(0xEB), 0xD9] // U+6CC6 <cjk>
	`泔`: [u8(0xEB), 0xDA] // U+6CD4 <cjk>
	`泠`: [u8(0xEB), 0xDB] // U+6CE0 <cjk>
	`泫`: [u8(0xEB), 0xDC] // U+6CEB <cjk>
	`泮`: [u8(0xEB), 0xDD] // U+6CEE <cjk>
	`𣳾`: [u8(0xEB), 0xDE] // U+23CFE <cjk>
	`洄`: [u8(0xEB), 0xDF] // U+6D04 <cjk>
	`洎`: [u8(0xEB), 0xE0] // U+6D0E <cjk>
	`洮`: [u8(0xEB), 0xE1] // U+6D2E <cjk>
	`洱`: [u8(0xEB), 0xE2] // U+6D31 <cjk>
	`洹`: [u8(0xEB), 0xE3] // U+6D39 <cjk>
	`洿`: [u8(0xEB), 0xE4] // U+6D3F <cjk>
	`浘`: [u8(0xEB), 0xE5] // U+6D58 <cjk>
	`浥`: [u8(0xEB), 0xE6] // U+6D65 <cjk>
	`海`: [u8(0xEB), 0xE7] // U+FA45 CJK COMPATIBILITY IDEOGRAPH-FA45
	`涂`: [u8(0xEB), 0xE8] // U+6D82 <cjk>
	`涇`: [u8(0xEB), 0xE9] // U+6D87 <cjk>
	`涉`: [u8(0xEB), 0xEA] // U+6D89 <cjk>
	`涔`: [u8(0xEB), 0xEB] // U+6D94 <cjk>
	`涪`: [u8(0xEB), 0xEC] // U+6DAA <cjk>
	`涬`: [u8(0xEB), 0xED] // U+6DAC <cjk>
	`涿`: [u8(0xEB), 0xEE] // U+6DBF <cjk>
	`淄`: [u8(0xEB), 0xEF] // U+6DC4 <cjk>
	`淖`: [u8(0xEB), 0xF0] // U+6DD6 <cjk>
	`淚`: [u8(0xEB), 0xF1] // U+6DDA <cjk>
	`淛`: [u8(0xEB), 0xF2] // U+6DDB <cjk>
	`淝`: [u8(0xEB), 0xF3] // U+6DDD <cjk>
	`淼`: [u8(0xEB), 0xF4] // U+6DFC <cjk>
	`渚`: [u8(0xEB), 0xF5] // U+FA46 CJK COMPATIBILITY IDEOGRAPH-FA46
	`渴`: [u8(0xEB), 0xF6] // U+6E34 <cjk>
	`湄`: [u8(0xEB), 0xF7] // U+6E44 <cjk>
	`湜`: [u8(0xEB), 0xF8] // U+6E5C <cjk>
	`湞`: [u8(0xEB), 0xF9] // U+6E5E <cjk>
	`溫`: [u8(0xEB), 0xFA] // U+6EAB <cjk>
	`溱`: [u8(0xEB), 0xFB] // U+6EB1 <cjk>
	`滁`: [u8(0xEB), 0xFC] // U+6EC1 <cjk>
	`滇`: [u8(0xEC), 0x40] // U+6EC7 <cjk>
	`滎`: [u8(0xEC), 0x41] // U+6ECE <cjk>
	`漐`: [u8(0xEC), 0x42] // U+6F10 <cjk>
	`漚`: [u8(0xEC), 0x43] // U+6F1A <cjk>
	`漢`: [u8(0xEC), 0x44] // U+FA47 CJK COMPATIBILITY IDEOGRAPH-FA47
	`漪`: [u8(0xEC), 0x45] // U+6F2A <cjk>
	`漯`: [u8(0xEC), 0x46] // U+6F2F <cjk>
	`漳`: [u8(0xEC), 0x47] // U+6F33 <cjk>
	`潑`: [u8(0xEC), 0x48] // U+6F51 <cjk>
	`潙`: [u8(0xEC), 0x49] // U+6F59 <cjk>
	`潞`: [u8(0xEC), 0x4A] // U+6F5E <cjk>
	`潡`: [u8(0xEC), 0x4B] // U+6F61 <cjk>
	`潢`: [u8(0xEC), 0x4C] // U+6F62 <cjk>
	`潾`: [u8(0xEC), 0x4D] // U+6F7E <cjk>
	`澈`: [u8(0xEC), 0x4E] // U+6F88 <cjk>
	`澌`: [u8(0xEC), 0x4F] // U+6F8C <cjk>
	`澍`: [u8(0xEC), 0x50] // U+6F8D <cjk>
	`澔`: [u8(0xEC), 0x51] // U+6F94 <cjk>
	`澠`: [u8(0xEC), 0x52] // U+6FA0 <cjk>
	`澧`: [u8(0xEC), 0x53] // U+6FA7 <cjk>
	`澶`: [u8(0xEC), 0x54] // U+6FB6 <cjk>
	`澼`: [u8(0xEC), 0x55] // U+6FBC <cjk>
	`濇`: [u8(0xEC), 0x56] // U+6FC7 <cjk>
	`濊`: [u8(0xEC), 0x57] // U+6FCA <cjk>
	`濹`: [u8(0xEC), 0x58] // U+6FF9 <cjk>
	`濰`: [u8(0xEC), 0x59] // U+6FF0 <cjk>
	`濵`: [u8(0xEC), 0x5A] // U+6FF5 <cjk>
	`瀅`: [u8(0xEC), 0x5B] // U+7005 <cjk>
	`瀆`: [u8(0xEC), 0x5C] // U+7006 <cjk>
	`瀨`: [u8(0xEC), 0x5D] // U+7028 <cjk>
	`灊`: [u8(0xEC), 0x5E] // U+704A <cjk>
	`灝`: [u8(0xEC), 0x5F] // U+705D <cjk>
	`灞`: [u8(0xEC), 0x60] // U+705E <cjk>
	`灎`: [u8(0xEC), 0x61] // U+704E <cjk>
	`灤`: [u8(0xEC), 0x62] // U+7064 <cjk>
	`灵`: [u8(0xEC), 0x63] // U+7075 <cjk>
	`炅`: [u8(0xEC), 0x64] // U+7085 <cjk>
	`炤`: [u8(0xEC), 0x65] // U+70A4 <cjk>
	`炫`: [u8(0xEC), 0x66] // U+70AB <cjk>
	`炷`: [u8(0xEC), 0x67] // U+70B7 <cjk>
	`烔`: [u8(0xEC), 0x68] // U+70D4 <cjk>
	`烘`: [u8(0xEC), 0x69] // U+70D8 <cjk>
	`烤`: [u8(0xEC), 0x6A] // U+70E4 <cjk>
	`焏`: [u8(0xEC), 0x6B] // U+710F <cjk>
	`焫`: [u8(0xEC), 0x6C] // U+712B <cjk>
	`焞`: [u8(0xEC), 0x6D] // U+711E <cjk>
	`焠`: [u8(0xEC), 0x6E] // U+7120 <cjk>
	`焮`: [u8(0xEC), 0x6F] // U+712E <cjk>
	`焰`: [u8(0xEC), 0x70] // U+7130 <cjk>
	`煆`: [u8(0xEC), 0x71] // U+7146 <cjk>
	`煇`: [u8(0xEC), 0x72] // U+7147 <cjk>
	`煑`: [u8(0xEC), 0x73] // U+7151 <cjk>
	`煮`: [u8(0xEC), 0x74] // U+FA48 CJK COMPATIBILITY IDEOGRAPH-FA48
	`煒`: [u8(0xEC), 0x75] // U+7152 <cjk>
	`煜`: [u8(0xEC), 0x76] // U+715C <cjk>
	`煠`: [u8(0xEC), 0x77] // U+7160 <cjk>
	`煨`: [u8(0xEC), 0x78] // U+7168 <cjk>
	`凞`: [u8(0xEC), 0x79] // U+FA15 CJK COMPATIBILITY IDEOGRAPH-FA15
	`熅`: [u8(0xEC), 0x7A] // U+7185 <cjk>
	`熇`: [u8(0xEC), 0x7B] // U+7187 <cjk>
	`熒`: [u8(0xEC), 0x7C] // U+7192 <cjk>
	`燁`: [u8(0xEC), 0x7D] // U+71C1 <cjk>
	`熺`: [u8(0xEC), 0x7E] // U+71BA <cjk>
	`燄`: [u8(0xEC), 0x80] // U+71C4 <cjk>
	`燾`: [u8(0xEC), 0x81] // U+71FE <cjk>
	`爀`: [u8(0xEC), 0x82] // U+7200 <cjk>
	`爕`: [u8(0xEC), 0x83] // U+7215 <cjk>
	`牕`: [u8(0xEC), 0x84] // U+7255 <cjk>
	`牖`: [u8(0xEC), 0x85] // U+7256 <cjk>
	`㸿`: [u8(0xEC), 0x86] // U+3E3F <cjk>
	`犍`: [u8(0xEC), 0x87] // U+728D <cjk>
	`犛`: [u8(0xEC), 0x88] // U+729B <cjk>
	`犾`: [u8(0xEC), 0x89] // U+72BE <cjk>
	`狀`: [u8(0xEC), 0x8A] // U+72C0 <cjk>
	`狻`: [u8(0xEC), 0x8B] // U+72FB <cjk>
	`𤟱`: [u8(0xEC), 0x8C] // U+247F1 <cjk>
	`猧`: [u8(0xEC), 0x8D] // U+7327 <cjk>
	`猨`: [u8(0xEC), 0x8E] // U+7328 <cjk>
	`猪`: [u8(0xEC), 0x8F] // U+FA16 CJK COMPATIBILITY IDEOGRAPH-FA16
	`獐`: [u8(0xEC), 0x90] // U+7350 <cjk>
	`獦`: [u8(0xEC), 0x91] // U+7366 <cjk>
	`獼`: [u8(0xEC), 0x92] // U+737C <cjk>
	`玕`: [u8(0xEC), 0x93] // U+7395 <cjk>
	`玟`: [u8(0xEC), 0x94] // U+739F <cjk>
	`玠`: [u8(0xEC), 0x95] // U+73A0 <cjk>
	`玢`: [u8(0xEC), 0x96] // U+73A2 <cjk>
	`玦`: [u8(0xEC), 0x97] // U+73A6 <cjk>
	`玫`: [u8(0xEC), 0x98] // U+73AB <cjk>
	`珉`: [u8(0xEC), 0x99] // U+73C9 <cjk>
	`珏`: [u8(0xEC), 0x9A] // U+73CF <cjk>
	`珖`: [u8(0xEC), 0x9B] // U+73D6 <cjk>
	`珙`: [u8(0xEC), 0x9C] // U+73D9 <cjk>
	`珣`: [u8(0xEC), 0x9D] // U+73E3 <cjk>
	`珩`: [u8(0xEC), 0x9E] // U+73E9 <cjk>
	`琇`: [u8(0xEC), 0x9F] // U+7407 <cjk>
	`琊`: [u8(0xEC), 0xA0] // U+740A <cjk>
	`琚`: [u8(0xEC), 0xA1] // U+741A <cjk>
	`琛`: [u8(0xEC), 0xA2] // U+741B <cjk>
	`琢`: [u8(0xEC), 0xA3] // U+FA4A CJK COMPATIBILITY IDEOGRAPH-FA4A
	`琦`: [u8(0xEC), 0xA4] // U+7426 <cjk>
	`琨`: [u8(0xEC), 0xA5] // U+7428 <cjk>
	`琪`: [u8(0xEC), 0xA6] // U+742A <cjk>
	`琫`: [u8(0xEC), 0xA7] // U+742B <cjk>
	`琬`: [u8(0xEC), 0xA8] // U+742C <cjk>
	`琮`: [u8(0xEC), 0xA9] // U+742E <cjk>
	`琯`: [u8(0xEC), 0xAA] // U+742F <cjk>
	`琰`: [u8(0xEC), 0xAB] // U+7430 <cjk>
	`瑄`: [u8(0xEC), 0xAC] // U+7444 <cjk>
	`瑆`: [u8(0xEC), 0xAD] // U+7446 <cjk>
	`瑇`: [u8(0xEC), 0xAE] // U+7447 <cjk>
	`瑋`: [u8(0xEC), 0xAF] // U+744B <cjk>
	`瑗`: [u8(0xEC), 0xB0] // U+7457 <cjk>
	`瑢`: [u8(0xEC), 0xB1] // U+7462 <cjk>
	`瑫`: [u8(0xEC), 0xB2] // U+746B <cjk>
	`瑭`: [u8(0xEC), 0xB3] // U+746D <cjk>
	`璆`: [u8(0xEC), 0xB4] // U+7486 <cjk>
	`璇`: [u8(0xEC), 0xB5] // U+7487 <cjk>
	`璉`: [u8(0xEC), 0xB6] // U+7489 <cjk>
	`璘`: [u8(0xEC), 0xB7] // U+7498 <cjk>
	`璜`: [u8(0xEC), 0xB8] // U+749C <cjk>
	`璟`: [u8(0xEC), 0xB9] // U+749F <cjk>
	`璣`: [u8(0xEC), 0xBA] // U+74A3 <cjk>
	`璐`: [u8(0xEC), 0xBB] // U+7490 <cjk>
	`璦`: [u8(0xEC), 0xBC] // U+74A6 <cjk>
	`璨`: [u8(0xEC), 0xBD] // U+74A8 <cjk>
	`璩`: [u8(0xEC), 0xBE] // U+74A9 <cjk>
	`璵`: [u8(0xEC), 0xBF] // U+74B5 <cjk>
	`璿`: [u8(0xEC), 0xC0] // U+74BF <cjk>
	`瓈`: [u8(0xEC), 0xC1] // U+74C8 <cjk>
	`瓉`: [u8(0xEC), 0xC2] // U+74C9 <cjk>
	`瓚`: [u8(0xEC), 0xC3] // U+74DA <cjk>
	`瓿`: [u8(0xEC), 0xC4] // U+74FF <cjk>
	`甁`: [u8(0xEC), 0xC5] // U+7501 <cjk>
	`甗`: [u8(0xEC), 0xC6] // U+7517 <cjk>
	`甯`: [u8(0xEC), 0xC7] // U+752F <cjk>
	`畯`: [u8(0xEC), 0xC8] // U+756F <cjk>
	`畹`: [u8(0xEC), 0xC9] // U+7579 <cjk>
	`疒`: [u8(0xEC), 0xCA] // U+7592 <cjk>
	`㽲`: [u8(0xEC), 0xCB] // U+3F72 <cjk>
	`痎`: [u8(0xEC), 0xCC] // U+75CE <cjk>
	`痤`: [u8(0xEC), 0xCD] // U+75E4 <cjk>
	`瘀`: [u8(0xEC), 0xCE] // U+7600 <cjk>
	`瘂`: [u8(0xEC), 0xCF] // U+7602 <cjk>
	`瘈`: [u8(0xEC), 0xD0] // U+7608 <cjk>
	`瘕`: [u8(0xEC), 0xD1] // U+7615 <cjk>
	`瘖`: [u8(0xEC), 0xD2] // U+7616 <cjk>
	`瘙`: [u8(0xEC), 0xD3] // U+7619 <cjk>
	`瘞`: [u8(0xEC), 0xD4] // U+761E <cjk>
	`瘭`: [u8(0xEC), 0xD5] // U+762D <cjk>
	`瘵`: [u8(0xEC), 0xD6] // U+7635 <cjk>
	`癃`: [u8(0xEC), 0xD7] // U+7643 <cjk>
	`癋`: [u8(0xEC), 0xD8] // U+764B <cjk>
	`癤`: [u8(0xEC), 0xD9] // U+7664 <cjk>
	`癥`: [u8(0xEC), 0xDA] // U+7665 <cjk>
	`癭`: [u8(0xEC), 0xDB] // U+766D <cjk>
	`癯`: [u8(0xEC), 0xDC] // U+766F <cjk>
	`癱`: [u8(0xEC), 0xDD] // U+7671 <cjk>
	`皁`: [u8(0xEC), 0xDE] // U+7681 <cjk>
	`皛`: [u8(0xEC), 0xDF] // U+769B <cjk>
	`皝`: [u8(0xEC), 0xE0] // U+769D <cjk>
	`皞`: [u8(0xEC), 0xE1] // U+769E <cjk>
	`皦`: [u8(0xEC), 0xE2] // U+76A6 <cjk>
	`皪`: [u8(0xEC), 0xE3] // U+76AA <cjk>
	`皶`: [u8(0xEC), 0xE4] // U+76B6 <cjk>
	`盅`: [u8(0xEC), 0xE5] // U+76C5 <cjk>
	`盌`: [u8(0xEC), 0xE6] // U+76CC <cjk>
	`盎`: [u8(0xEC), 0xE7] // U+76CE <cjk>
	`盔`: [u8(0xEC), 0xE8] // U+76D4 <cjk>
	`盦`: [u8(0xEC), 0xE9] // U+76E6 <cjk>
	`盱`: [u8(0xEC), 0xEA] // U+76F1 <cjk>
	`盼`: [u8(0xEC), 0xEB] // U+76FC <cjk>
	`眊`: [u8(0xEC), 0xEC] // U+770A <cjk>
	`眙`: [u8(0xEC), 0xED] // U+7719 <cjk>
	`眴`: [u8(0xEC), 0xEE] // U+7734 <cjk>
	`眶`: [u8(0xEC), 0xEF] // U+7736 <cjk>
	`睆`: [u8(0xEC), 0xF0] // U+7746 <cjk>
	`睍`: [u8(0xEC), 0xF1] // U+774D <cjk>
	`睎`: [u8(0xEC), 0xF2] // U+774E <cjk>
	`睜`: [u8(0xEC), 0xF3] // U+775C <cjk>
	`睟`: [u8(0xEC), 0xF4] // U+775F <cjk>
	`睢`: [u8(0xEC), 0xF5] // U+7762 <cjk>
	`睺`: [u8(0xEC), 0xF6] // U+777A <cjk>
	`瞀`: [u8(0xEC), 0xF7] // U+7780 <cjk>
	`瞔`: [u8(0xEC), 0xF8] // U+7794 <cjk>
	`瞪`: [u8(0xEC), 0xF9] // U+77AA <cjk>
	`矠`: [u8(0xEC), 0xFA] // U+77E0 <cjk>
	`砭`: [u8(0xEC), 0xFB] // U+782D <cjk>
	`𥒎`: [u8(0xEC), 0xFC] // U+2548E <cjk>
	`硃`: [u8(0xED), 0x40] // U+7843 <cjk>
	`硎`: [u8(0xED), 0x41] // U+784E <cjk>
	`硏`: [u8(0xED), 0x42] // U+784F <cjk>
	`硑`: [u8(0xED), 0x43] // U+7851 <cjk>
	`硨`: [u8(0xED), 0x44] // U+7868 <cjk>
	`确`: [u8(0xED), 0x45] // U+786E <cjk>
	`碑`: [u8(0xED), 0x46] // U+FA4B CJK COMPATIBILITY IDEOGRAPH-FA4B
	`碰`: [u8(0xED), 0x47] // U+78B0 <cjk>
	`𥔎`: [u8(0xED), 0x48] // U+2550E <cjk>
	`碭`: [u8(0xED), 0x49] // U+78AD <cjk>
	`磤`: [u8(0xED), 0x4A] // U+78E4 <cjk>
	`磲`: [u8(0xED), 0x4B] // U+78F2 <cjk>
	`礀`: [u8(0xED), 0x4C] // U+7900 <cjk>
	`磷`: [u8(0xED), 0x4D] // U+78F7 <cjk>
	`礜`: [u8(0xED), 0x4E] // U+791C <cjk>
	`礮`: [u8(0xED), 0x4F] // U+792E <cjk>
	`礱`: [u8(0xED), 0x50] // U+7931 <cjk>
	`礴`: [u8(0xED), 0x51] // U+7934 <cjk>
	`社`: [u8(0xED), 0x52] // U+FA4C CJK COMPATIBILITY IDEOGRAPH-FA4C
	`祉`: [u8(0xED), 0x53] // U+FA4D CJK COMPATIBILITY IDEOGRAPH-FA4D
	`祅`: [u8(0xED), 0x54] // U+7945 <cjk>
	`祆`: [u8(0xED), 0x55] // U+7946 <cjk>
	`祈`: [u8(0xED), 0x56] // U+FA4E CJK COMPATIBILITY IDEOGRAPH-FA4E
	`祐`: [u8(0xED), 0x57] // U+FA4F CJK COMPATIBILITY IDEOGRAPH-FA4F
	`祖`: [u8(0xED), 0x58] // U+FA50 CJK COMPATIBILITY IDEOGRAPH-FA50
	`祜`: [u8(0xED), 0x59] // U+795C <cjk>
	`祝`: [u8(0xED), 0x5A] // U+FA51 CJK COMPATIBILITY IDEOGRAPH-FA51
	`神`: [u8(0xED), 0x5B] // U+FA19 CJK COMPATIBILITY IDEOGRAPH-FA19
	`祥`: [u8(0xED), 0x5C] // U+FA1A CJK COMPATIBILITY IDEOGRAPH-FA1A
	`祹`: [u8(0xED), 0x5D] // U+7979 <cjk>
	`禍`: [u8(0xED), 0x5E] // U+FA52 CJK COMPATIBILITY IDEOGRAPH-FA52
	`禎`: [u8(0xED), 0x5F] // U+FA53 CJK COMPATIBILITY IDEOGRAPH-FA53
	`福`: [u8(0xED), 0x60] // U+FA1B CJK COMPATIBILITY IDEOGRAPH-FA1B
	`禘`: [u8(0xED), 0x61] // U+7998 <cjk>
	`禱`: [u8(0xED), 0x62] // U+79B1 <cjk>
	`禸`: [u8(0xED), 0x63] // U+79B8 <cjk>
	`秈`: [u8(0xED), 0x64] // U+79C8 <cjk>
	`秊`: [u8(0xED), 0x65] // U+79CA <cjk>
	`𥝱`: [u8(0xED), 0x66] // U+25771 <cjk>
	`秔`: [u8(0xED), 0x67] // U+79D4 <cjk>
	`秞`: [u8(0xED), 0x68] // U+79DE <cjk>
	`秫`: [u8(0xED), 0x69] // U+79EB <cjk>
	`秭`: [u8(0xED), 0x6A] // U+79ED <cjk>
	`稃`: [u8(0xED), 0x6B] // U+7A03 <cjk>
	`穀`: [u8(0xED), 0x6C] // U+FA54 CJK COMPATIBILITY IDEOGRAPH-FA54
	`稹`: [u8(0xED), 0x6D] // U+7A39 <cjk>
	`穝`: [u8(0xED), 0x6E] // U+7A5D <cjk>
	`穭`: [u8(0xED), 0x6F] // U+7A6D <cjk>
	`突`: [u8(0xED), 0x70] // U+FA55 CJK COMPATIBILITY IDEOGRAPH-FA55
	`窅`: [u8(0xED), 0x71] // U+7A85 <cjk>
	`窠`: [u8(0xED), 0x72] // U+7AA0 <cjk>
	`𥧄`: [u8(0xED), 0x73] // U+259C4 <cjk>
	`窳`: [u8(0xED), 0x74] // U+7AB3 <cjk>
	`窻`: [u8(0xED), 0x75] // U+7ABB <cjk>
	`竎`: [u8(0xED), 0x76] // U+7ACE <cjk>
	`竫`: [u8(0xED), 0x77] // U+7AEB <cjk>
	`竽`: [u8(0xED), 0x78] // U+7AFD <cjk>
	`笒`: [u8(0xED), 0x79] // U+7B12 <cjk>
	`笭`: [u8(0xED), 0x7A] // U+7B2D <cjk>
	`笻`: [u8(0xED), 0x7B] // U+7B3B <cjk>
	`筇`: [u8(0xED), 0x7C] // U+7B47 <cjk>
	`筎`: [u8(0xED), 0x7D] // U+7B4E <cjk>
	`筠`: [u8(0xED), 0x7E] // U+7B60 <cjk>
	`筭`: [u8(0xED), 0x80] // U+7B6D <cjk>
	`筯`: [u8(0xED), 0x81] // U+7B6F <cjk>
	`筲`: [u8(0xED), 0x82] // U+7B72 <cjk>
	`箞`: [u8(0xED), 0x83] // U+7B9E <cjk>
	`節`: [u8(0xED), 0x84] // U+FA56 CJK COMPATIBILITY IDEOGRAPH-FA56
	`篗`: [u8(0xED), 0x85] // U+7BD7 <cjk>
	`篙`: [u8(0xED), 0x86] // U+7BD9 <cjk>
	`簁`: [u8(0xED), 0x87] // U+7C01 <cjk>
	`簱`: [u8(0xED), 0x88] // U+7C31 <cjk>
	`簞`: [u8(0xED), 0x89] // U+7C1E <cjk>
	`簠`: [u8(0xED), 0x8A] // U+7C20 <cjk>
	`簳`: [u8(0xED), 0x8B] // U+7C33 <cjk>
	`簶`: [u8(0xED), 0x8C] // U+7C36 <cjk>
	`䉤`: [u8(0xED), 0x8D] // U+4264 <cjk>
	`𥶡`: [u8(0xED), 0x8E] // U+25DA1 <cjk>
	`籙`: [u8(0xED), 0x8F] // U+7C59 <cjk>
	`籭`: [u8(0xED), 0x90] // U+7C6D <cjk>
	`籹`: [u8(0xED), 0x91] // U+7C79 <cjk>
	`粏`: [u8(0xED), 0x92] // U+7C8F <cjk>
	`粔`: [u8(0xED), 0x93] // U+7C94 <cjk>
	`粠`: [u8(0xED), 0x94] // U+7CA0 <cjk>
	`粼`: [u8(0xED), 0x95] // U+7CBC <cjk>
	`糕`: [u8(0xED), 0x96] // U+7CD5 <cjk>
	`糙`: [u8(0xED), 0x97] // U+7CD9 <cjk>
	`糝`: [u8(0xED), 0x98] // U+7CDD <cjk>
	`紇`: [u8(0xED), 0x99] // U+7D07 <cjk>
	`紈`: [u8(0xED), 0x9A] // U+7D08 <cjk>
	`紓`: [u8(0xED), 0x9B] // U+7D13 <cjk>
	`紝`: [u8(0xED), 0x9C] // U+7D1D <cjk>
	`紣`: [u8(0xED), 0x9D] // U+7D23 <cjk>
	`紱`: [u8(0xED), 0x9E] // U+7D31 <cjk>
	`絁`: [u8(0xED), 0x9F] // U+7D41 <cjk>
	`絈`: [u8(0xED), 0xA0] // U+7D48 <cjk>
	`絓`: [u8(0xED), 0xA1] // U+7D53 <cjk>
	`絜`: [u8(0xED), 0xA2] // U+7D5C <cjk>
	`絺`: [u8(0xED), 0xA3] // U+7D7A <cjk>
	`綃`: [u8(0xED), 0xA4] // U+7D83 <cjk>
	`綋`: [u8(0xED), 0xA5] // U+7D8B <cjk>
	`綠`: [u8(0xED), 0xA6] // U+7DA0 <cjk>
	`綦`: [u8(0xED), 0xA7] // U+7DA6 <cjk>
	`緂`: [u8(0xED), 0xA8] // U+7DC2 <cjk>
	`緌`: [u8(0xED), 0xA9] // U+7DCC <cjk>
	`緖`: [u8(0xED), 0xAA] // U+7DD6 <cjk>
	`緣`: [u8(0xED), 0xAB] // U+7DE3 <cjk>
	`練`: [u8(0xED), 0xAC] // U+FA57 CJK COMPATIBILITY IDEOGRAPH-FA57
	`縨`: [u8(0xED), 0xAD] // U+7E28 <cjk>
	`縈`: [u8(0xED), 0xAE] // U+7E08 <cjk>
	`縑`: [u8(0xED), 0xAF] // U+7E11 <cjk>
	`縕`: [u8(0xED), 0xB0] // U+7E15 <cjk>
	`繁`: [u8(0xED), 0xB1] // U+FA59 CJK COMPATIBILITY IDEOGRAPH-FA59
	`繇`: [u8(0xED), 0xB2] // U+7E47 <cjk>
	`繒`: [u8(0xED), 0xB3] // U+7E52 <cjk>
	`繡`: [u8(0xED), 0xB4] // U+7E61 <cjk>
	`纊`: [u8(0xED), 0xB5] // U+7E8A <cjk>
	`纍`: [u8(0xED), 0xB6] // U+7E8D <cjk>
	`罇`: [u8(0xED), 0xB7] // U+7F47 <cjk>
	`署`: [u8(0xED), 0xB8] // U+FA5A CJK COMPATIBILITY IDEOGRAPH-FA5A
	`羑`: [u8(0xED), 0xB9] // U+7F91 <cjk>
	`羗`: [u8(0xED), 0xBA] // U+7F97 <cjk>
	`羿`: [u8(0xED), 0xBB] // U+7FBF <cjk>
	`翎`: [u8(0xED), 0xBC] // U+7FCE <cjk>
	`翛`: [u8(0xED), 0xBD] // U+7FDB <cjk>
	`翟`: [u8(0xED), 0xBE] // U+7FDF <cjk>
	`翬`: [u8(0xED), 0xBF] // U+7FEC <cjk>
	`翮`: [u8(0xED), 0xC0] // U+7FEE <cjk>
	`翺`: [u8(0xED), 0xC1] // U+7FFA <cjk>
	`者`: [u8(0xED), 0xC2] // U+FA5B CJK COMPATIBILITY IDEOGRAPH-FA5B
	`耔`: [u8(0xED), 0xC3] // U+8014 <cjk>
	`耦`: [u8(0xED), 0xC4] // U+8026 <cjk>
	`耵`: [u8(0xED), 0xC5] // U+8035 <cjk>
	`耷`: [u8(0xED), 0xC6] // U+8037 <cjk>
	`耼`: [u8(0xED), 0xC7] // U+803C <cjk>
	`胊`: [u8(0xED), 0xC8] // U+80CA <cjk>
	`胗`: [u8(0xED), 0xC9] // U+80D7 <cjk>
	`胠`: [u8(0xED), 0xCA] // U+80E0 <cjk>
	`胳`: [u8(0xED), 0xCB] // U+80F3 <cjk>
	`脘`: [u8(0xED), 0xCC] // U+8118 <cjk>
	`腊`: [u8(0xED), 0xCD] // U+814A <cjk>
	`腠`: [u8(0xED), 0xCE] // U+8160 <cjk>
	`腧`: [u8(0xED), 0xCF] // U+8167 <cjk>
	`腨`: [u8(0xED), 0xD0] // U+8168 <cjk>
	`腭`: [u8(0xED), 0xD1] // U+816D <cjk>
	`膻`: [u8(0xED), 0xD2] // U+81BB <cjk>
	`臊`: [u8(0xED), 0xD3] // U+81CA <cjk>
	`臏`: [u8(0xED), 0xD4] // U+81CF <cjk>
	`臗`: [u8(0xED), 0xD5] // U+81D7 <cjk>
	`臭`: [u8(0xED), 0xD6] // U+FA5C CJK COMPATIBILITY IDEOGRAPH-FA5C
	`䑓`: [u8(0xED), 0xD7] // U+4453 <cjk>
	`䑛`: [u8(0xED), 0xD8] // U+445B <cjk>
	`艠`: [u8(0xED), 0xD9] // U+8260 <cjk>
	`艴`: [u8(0xED), 0xDA] // U+8274 <cjk>
	`𦫿`: [u8(0xED), 0xDB] // U+26AFF <cjk>
	`芎`: [u8(0xED), 0xDC] // U+828E <cjk>
	`芡`: [u8(0xED), 0xDD] // U+82A1 <cjk>
	`芣`: [u8(0xED), 0xDE] // U+82A3 <cjk>
	`芤`: [u8(0xED), 0xDF] // U+82A4 <cjk>
	`芩`: [u8(0xED), 0xE0] // U+82A9 <cjk>
	`芮`: [u8(0xED), 0xE1] // U+82AE <cjk>
	`芷`: [u8(0xED), 0xE2] // U+82B7 <cjk>
	`芾`: [u8(0xED), 0xE3] // U+82BE <cjk>
	`芿`: [u8(0xED), 0xE4] // U+82BF <cjk>
	`苆`: [u8(0xED), 0xE5] // U+82C6 <cjk>
	`苕`: [u8(0xED), 0xE6] // U+82D5 <cjk>
	`苽`: [u8(0xED), 0xE7] // U+82FD <cjk>
	`苾`: [u8(0xED), 0xE8] // U+82FE <cjk>
	`茀`: [u8(0xED), 0xE9] // U+8300 <cjk>
	`茁`: [u8(0xED), 0xEA] // U+8301 <cjk>
	`荢`: [u8(0xED), 0xEB] // U+8362 <cjk>
	`茢`: [u8(0xED), 0xEC] // U+8322 <cjk>
	`茭`: [u8(0xED), 0xED] // U+832D <cjk>
	`茺`: [u8(0xED), 0xEE] // U+833A <cjk>
	`荃`: [u8(0xED), 0xEF] // U+8343 <cjk>
	`荇`: [u8(0xED), 0xF0] // U+8347 <cjk>
	`荑`: [u8(0xED), 0xF1] // U+8351 <cjk>
	`荕`: [u8(0xED), 0xF2] // U+8355 <cjk>
	`荽`: [u8(0xED), 0xF3] // U+837D <cjk>
	`莆`: [u8(0xED), 0xF4] // U+8386 <cjk>
	`莒`: [u8(0xED), 0xF5] // U+8392 <cjk>
	`莘`: [u8(0xED), 0xF6] // U+8398 <cjk>
	`莧`: [u8(0xED), 0xF7] // U+83A7 <cjk>
	`莩`: [u8(0xED), 0xF8] // U+83A9 <cjk>
	`莿`: [u8(0xED), 0xF9] // U+83BF <cjk>
	`菀`: [u8(0xED), 0xFA] // U+83C0 <cjk>
	`菇`: [u8(0xED), 0xFB] // U+83C7 <cjk>
	`菏`: [u8(0xED), 0xFC] // U+83CF <cjk>
	`菑`: [u8(0xEE), 0x40] // U+83D1 <cjk>
	`菡`: [u8(0xEE), 0x41] // U+83E1 <cjk>
	`菪`: [u8(0xEE), 0x42] // U+83EA <cjk>
	`萁`: [u8(0xEE), 0x43] // U+8401 <cjk>
	`萆`: [u8(0xEE), 0x44] // U+8406 <cjk>
	`萊`: [u8(0xEE), 0x45] // U+840A <cjk>
	`著`: [u8(0xEE), 0x46] // U+FA5F CJK COMPATIBILITY IDEOGRAPH-FA5F
	`葈`: [u8(0xEE), 0x47] // U+8448 <cjk>
	`葟`: [u8(0xEE), 0x48] // U+845F <cjk>
	`葰`: [u8(0xEE), 0x49] // U+8470 <cjk>
	`葳`: [u8(0xEE), 0x4A] // U+8473 <cjk>
	`蒅`: [u8(0xEE), 0x4B] // U+8485 <cjk>
	`蒞`: [u8(0xEE), 0x4C] // U+849E <cjk>
	`蒯`: [u8(0xEE), 0x4D] // U+84AF <cjk>
	`蒴`: [u8(0xEE), 0x4E] // U+84B4 <cjk>
	`蒺`: [u8(0xEE), 0x4F] // U+84BA <cjk>
	`蓀`: [u8(0xEE), 0x50] // U+84C0 <cjk>
	`蓂`: [u8(0xEE), 0x51] // U+84C2 <cjk>
	`𦹀`: [u8(0xEE), 0x52] // U+26E40 <cjk>
	`蔲`: [u8(0xEE), 0x53] // U+8532 <cjk>
	`蔞`: [u8(0xEE), 0x54] // U+851E <cjk>
	`蔣`: [u8(0xEE), 0x55] // U+8523 <cjk>
	`蔯`: [u8(0xEE), 0x56] // U+852F <cjk>
	`蕙`: [u8(0xEE), 0x57] // U+8559 <cjk>
	`蕤`: [u8(0xEE), 0x58] // U+8564 <cjk>
	`﨟`: [u8(0xEE), 0x59] // U+FA1F CJK COMPATIBILITY IDEOGRAPH-FA1F
	`薭`: [u8(0xEE), 0x5A] // U+85AD <cjk>
	`蕺`: [u8(0xEE), 0x5B] // U+857A <cjk>
	`薌`: [u8(0xEE), 0x5C] // U+858C <cjk>
	`薏`: [u8(0xEE), 0x5D] // U+858F <cjk>
	`薢`: [u8(0xEE), 0x5E] // U+85A2 <cjk>
	`薰`: [u8(0xEE), 0x5F] // U+85B0 <cjk>
	`藋`: [u8(0xEE), 0x60] // U+85CB <cjk>
	`藎`: [u8(0xEE), 0x61] // U+85CE <cjk>
	`藭`: [u8(0xEE), 0x62] // U+85ED <cjk>
	`蘒`: [u8(0xEE), 0x63] // U+8612 <cjk>
	`藿`: [u8(0xEE), 0x64] // U+85FF <cjk>
	`蘄`: [u8(0xEE), 0x65] // U+8604 <cjk>
	`蘅`: [u8(0xEE), 0x66] // U+8605 <cjk>
	`蘐`: [u8(0xEE), 0x67] // U+8610 <cjk>
	`𧃴`: [u8(0xEE), 0x68] // U+270F4 <cjk>
	`蘘`: [u8(0xEE), 0x69] // U+8618 <cjk>
	`蘩`: [u8(0xEE), 0x6A] // U+8629 <cjk>
	`蘸`: [u8(0xEE), 0x6B] // U+8638 <cjk>
	`虗`: [u8(0xEE), 0x6C] // U+8657 <cjk>
	`虛`: [u8(0xEE), 0x6D] // U+865B <cjk>
	`虜`: [u8(0xEE), 0x6E] // U+F936 CJK COMPATIBILITY IDEOGRAPH-F936
	`虢`: [u8(0xEE), 0x6F] // U+8662 <cjk>
	`䖝`: [u8(0xEE), 0x70] // U+459D <cjk>
	`虬`: [u8(0xEE), 0x71] // U+866C <cjk>
	`虵`: [u8(0xEE), 0x72] // U+8675 <cjk>
	`蚘`: [u8(0xEE), 0x73] // U+8698 <cjk>
	`蚸`: [u8(0xEE), 0x74] // U+86B8 <cjk>
	`蛺`: [u8(0xEE), 0x75] // U+86FA <cjk>
	`蛼`: [u8(0xEE), 0x76] // U+86FC <cjk>
	`蛽`: [u8(0xEE), 0x77] // U+86FD <cjk>
	`蜋`: [u8(0xEE), 0x78] // U+870B <cjk>
	`蝱`: [u8(0xEE), 0x79] // U+8771 <cjk>
	`螇`: [u8(0xEE), 0x7A] // U+8787 <cjk>
	`螈`: [u8(0xEE), 0x7B] // U+8788 <cjk>
	`螬`: [u8(0xEE), 0x7C] // U+87AC <cjk>
	`螭`: [u8(0xEE), 0x7D] // U+87AD <cjk>
	`螵`: [u8(0xEE), 0x7E] // U+87B5 <cjk>
	`䗪`: [u8(0xEE), 0x80] // U+45EA <cjk>
	`蟖`: [u8(0xEE), 0x81] // U+87D6 <cjk>
	`蟬`: [u8(0xEE), 0x82] // U+87EC <cjk>
	`蠆`: [u8(0xEE), 0x83] // U+8806 <cjk>
	`蠊`: [u8(0xEE), 0x84] // U+880A <cjk>
	`蠐`: [u8(0xEE), 0x85] // U+8810 <cjk>
	`蠔`: [u8(0xEE), 0x86] // U+8814 <cjk>
	`蠟`: [u8(0xEE), 0x87] // U+881F <cjk>
	`袘`: [u8(0xEE), 0x88] // U+8898 <cjk>
	`袪`: [u8(0xEE), 0x89] // U+88AA <cjk>
	`裊`: [u8(0xEE), 0x8A] // U+88CA <cjk>
	`裎`: [u8(0xEE), 0x8B] // U+88CE <cjk>
	`𧚄`: [u8(0xEE), 0x8C] // U+27684 <cjk>
	`裵`: [u8(0xEE), 0x8D] // U+88F5 <cjk>
	`褜`: [u8(0xEE), 0x8E] // U+891C <cjk>
	`褐`: [u8(0xEE), 0x8F] // U+FA60 CJK COMPATIBILITY IDEOGRAPH-FA60
	`褘`: [u8(0xEE), 0x90] // U+8918 <cjk>
	`褙`: [u8(0xEE), 0x91] // U+8919 <cjk>
	`褚`: [u8(0xEE), 0x92] // U+891A <cjk>
	`褧`: [u8(0xEE), 0x93] // U+8927 <cjk>
	`褰`: [u8(0xEE), 0x94] // U+8930 <cjk>
	`褲`: [u8(0xEE), 0x95] // U+8932 <cjk>
	`褹`: [u8(0xEE), 0x96] // U+8939 <cjk>
	`襀`: [u8(0xEE), 0x97] // U+8940 <cjk>
	`覔`: [u8(0xEE), 0x98] // U+8994 <cjk>
	`視`: [u8(0xEE), 0x99] // U+FA61 CJK COMPATIBILITY IDEOGRAPH-FA61
	`觔`: [u8(0xEE), 0x9A] // U+89D4 <cjk>
	`觥`: [u8(0xEE), 0x9B] // U+89E5 <cjk>
	`觶`: [u8(0xEE), 0x9C] // U+89F6 <cjk>
	`訒`: [u8(0xEE), 0x9D] // U+8A12 <cjk>
	`訕`: [u8(0xEE), 0x9E] // U+8A15 <cjk>
	`訢`: [u8(0xEE), 0x9F] // U+8A22 <cjk>
	`訷`: [u8(0xEE), 0xA0] // U+8A37 <cjk>
	`詇`: [u8(0xEE), 0xA1] // U+8A47 <cjk>
	`詎`: [u8(0xEE), 0xA2] // U+8A4E <cjk>
	`詝`: [u8(0xEE), 0xA3] // U+8A5D <cjk>
	`詡`: [u8(0xEE), 0xA4] // U+8A61 <cjk>
	`詵`: [u8(0xEE), 0xA5] // U+8A75 <cjk>
	`詹`: [u8(0xEE), 0xA6] // U+8A79 <cjk>
	`誧`: [u8(0xEE), 0xA7] // U+8AA7 <cjk>
	`諐`: [u8(0xEE), 0xA8] // U+8AD0 <cjk>
	`諟`: [u8(0xEE), 0xA9] // U+8ADF <cjk>
	`諴`: [u8(0xEE), 0xAA] // U+8AF4 <cjk>
	`諶`: [u8(0xEE), 0xAB] // U+8AF6 <cjk>
	`諸`: [u8(0xEE), 0xAC] // U+FA22 CJK COMPATIBILITY IDEOGRAPH-FA22
	`謁`: [u8(0xEE), 0xAD] // U+FA62 CJK COMPATIBILITY IDEOGRAPH-FA62
	`謹`: [u8(0xEE), 0xAE] // U+FA63 CJK COMPATIBILITY IDEOGRAPH-FA63
	`譆`: [u8(0xEE), 0xAF] // U+8B46 <cjk>
	`譔`: [u8(0xEE), 0xB0] // U+8B54 <cjk>
	`譙`: [u8(0xEE), 0xB1] // U+8B59 <cjk>
	`譩`: [u8(0xEE), 0xB2] // U+8B69 <cjk>
	`讝`: [u8(0xEE), 0xB3] // U+8B9D <cjk>
	`豉`: [u8(0xEE), 0xB4] // U+8C49 <cjk>
	`豨`: [u8(0xEE), 0xB5] // U+8C68 <cjk>
	`賓`: [u8(0xEE), 0xB6] // U+FA64 CJK COMPATIBILITY IDEOGRAPH-FA64
	`賡`: [u8(0xEE), 0xB7] // U+8CE1 <cjk>
	`賴`: [u8(0xEE), 0xB8] // U+8CF4 <cjk>
	`賸`: [u8(0xEE), 0xB9] // U+8CF8 <cjk>
	`賾`: [u8(0xEE), 0xBA] // U+8CFE <cjk>
	`贈`: [u8(0xEE), 0xBB] // U+FA65 CJK COMPATIBILITY IDEOGRAPH-FA65
	`贒`: [u8(0xEE), 0xBC] // U+8D12 <cjk>
	`贛`: [u8(0xEE), 0xBD] // U+8D1B <cjk>
	`趯`: [u8(0xEE), 0xBE] // U+8DAF <cjk>
	`跎`: [u8(0xEE), 0xBF] // U+8DCE <cjk>
	`跑`: [u8(0xEE), 0xC0] // U+8DD1 <cjk>
	`跗`: [u8(0xEE), 0xC1] // U+8DD7 <cjk>
	`踠`: [u8(0xEE), 0xC2] // U+8E20 <cjk>
	`踣`: [u8(0xEE), 0xC3] // U+8E23 <cjk>
	`踽`: [u8(0xEE), 0xC4] // U+8E3D <cjk>
	`蹰`: [u8(0xEE), 0xC5] // U+8E70 <cjk>
	`蹻`: [u8(0xEE), 0xC6] // U+8E7B <cjk>
	`𨉷`: [u8(0xEE), 0xC7] // U+28277 <cjk>
	`軀`: [u8(0xEE), 0xC8] // U+8EC0 <cjk>
	`䡄`: [u8(0xEE), 0xC9] // U+4844 <cjk>
	`軺`: [u8(0xEE), 0xCA] // U+8EFA <cjk>
	`輞`: [u8(0xEE), 0xCB] // U+8F1E <cjk>
	`輭`: [u8(0xEE), 0xCC] // U+8F2D <cjk>
	`輶`: [u8(0xEE), 0xCD] // U+8F36 <cjk>
	`轔`: [u8(0xEE), 0xCE] // U+8F54 <cjk>
	`𨏍`: [u8(0xEE), 0xCF] // U+283CD <cjk>
	`辦`: [u8(0xEE), 0xD0] // U+8FA6 <cjk>
	`辵`: [u8(0xEE), 0xD1] // U+8FB5 <cjk>
	`迤`: [u8(0xEE), 0xD2] // U+8FE4 <cjk>
	`迨`: [u8(0xEE), 0xD3] // U+8FE8 <cjk>
	`迮`: [u8(0xEE), 0xD4] // U+8FEE <cjk>
	`逈`: [u8(0xEE), 0xD5] // U+9008 <cjk>
	`逭`: [u8(0xEE), 0xD6] // U+902D <cjk>
	`逸`: [u8(0xEE), 0xD7] // U+FA67 CJK COMPATIBILITY IDEOGRAPH-FA67
	`邈`: [u8(0xEE), 0xD8] // U+9088 <cjk>
	`邕`: [u8(0xEE), 0xD9] // U+9095 <cjk>
	`邗`: [u8(0xEE), 0xDA] // U+9097 <cjk>
	`邙`: [u8(0xEE), 0xDB] // U+9099 <cjk>
	`邛`: [u8(0xEE), 0xDC] // U+909B <cjk>
	`邢`: [u8(0xEE), 0xDD] // U+90A2 <cjk>
	`邳`: [u8(0xEE), 0xDE] // U+90B3 <cjk>
	`邾`: [u8(0xEE), 0xDF] // U+90BE <cjk>
	`郄`: [u8(0xEE), 0xE0] // U+90C4 <cjk>
	`郅`: [u8(0xEE), 0xE1] // U+90C5 <cjk>
	`郇`: [u8(0xEE), 0xE2] // U+90C7 <cjk>
	`郗`: [u8(0xEE), 0xE3] // U+90D7 <cjk>
	`郝`: [u8(0xEE), 0xE4] // U+90DD <cjk>
	`郞`: [u8(0xEE), 0xE5] // U+90DE <cjk>
	`郯`: [u8(0xEE), 0xE6] // U+90EF <cjk>
	`郴`: [u8(0xEE), 0xE7] // U+90F4 <cjk>
	`都`: [u8(0xEE), 0xE8] // U+FA26 CJK COMPATIBILITY IDEOGRAPH-FA26
	`鄔`: [u8(0xEE), 0xE9] // U+9114 <cjk>
	`鄕`: [u8(0xEE), 0xEA] // U+9115 <cjk>
	`鄖`: [u8(0xEE), 0xEB] // U+9116 <cjk>
	`鄢`: [u8(0xEE), 0xEC] // U+9122 <cjk>
	`鄣`: [u8(0xEE), 0xED] // U+9123 <cjk>
	`鄧`: [u8(0xEE), 0xEE] // U+9127 <cjk>
	`鄯`: [u8(0xEE), 0xEF] // U+912F <cjk>
	`鄱`: [u8(0xEE), 0xF0] // U+9131 <cjk>
	`鄴`: [u8(0xEE), 0xF1] // U+9134 <cjk>
	`鄽`: [u8(0xEE), 0xF2] // U+913D <cjk>
	`酈`: [u8(0xEE), 0xF3] // U+9148 <cjk>
	`酛`: [u8(0xEE), 0xF4] // U+915B <cjk>
	`醃`: [u8(0xEE), 0xF5] // U+9183 <cjk>
	`醞`: [u8(0xEE), 0xF6] // U+919E <cjk>
	`醬`: [u8(0xEE), 0xF7] // U+91AC <cjk>
	`醱`: [u8(0xEE), 0xF8] // U+91B1 <cjk>
	`醼`: [u8(0xEE), 0xF9] // U+91BC <cjk>
	`釗`: [u8(0xEE), 0xFA] // U+91D7 <cjk>
	`釻`: [u8(0xEE), 0xFB] // U+91FB <cjk>
	`釤`: [u8(0xEE), 0xFC] // U+91E4 <cjk>
	`釥`: [u8(0xEF), 0x40] // U+91E5 <cjk>
	`釭`: [u8(0xEF), 0x41] // U+91ED <cjk>
	`釱`: [u8(0xEF), 0x42] // U+91F1 <cjk>
	`鈇`: [u8(0xEF), 0x43] // U+9207 <cjk>
	`鈐`: [u8(0xEF), 0x44] // U+9210 <cjk>
	`鈸`: [u8(0xEF), 0x45] // U+9238 <cjk>
	`鈹`: [u8(0xEF), 0x46] // U+9239 <cjk>
	`鈺`: [u8(0xEF), 0x47] // U+923A <cjk>
	`鈼`: [u8(0xEF), 0x48] // U+923C <cjk>
	`鉀`: [u8(0xEF), 0x49] // U+9240 <cjk>
	`鉃`: [u8(0xEF), 0x4A] // U+9243 <cjk>
	`鉏`: [u8(0xEF), 0x4B] // U+924F <cjk>
	`鉸`: [u8(0xEF), 0x4C] // U+9278 <cjk>
	`銈`: [u8(0xEF), 0x4D] // U+9288 <cjk>
	`鋂`: [u8(0xEF), 0x4E] // U+92C2 <cjk>
	`鋋`: [u8(0xEF), 0x4F] // U+92CB <cjk>
	`鋌`: [u8(0xEF), 0x50] // U+92CC <cjk>
	`鋓`: [u8(0xEF), 0x51] // U+92D3 <cjk>
	`鋠`: [u8(0xEF), 0x52] // U+92E0 <cjk>
	`鋿`: [u8(0xEF), 0x53] // U+92FF <cjk>
	`錄`: [u8(0xEF), 0x54] // U+9304 <cjk>
	`錟`: [u8(0xEF), 0x55] // U+931F <cjk>
	`錡`: [u8(0xEF), 0x56] // U+9321 <cjk>
	`錥`: [u8(0xEF), 0x57] // U+9325 <cjk>
	`鍈`: [u8(0xEF), 0x58] // U+9348 <cjk>
	`鍉`: [u8(0xEF), 0x59] // U+9349 <cjk>
	`鍊`: [u8(0xEF), 0x5A] // U+934A <cjk>
	`鍤`: [u8(0xEF), 0x5B] // U+9364 <cjk>
	`鍥`: [u8(0xEF), 0x5C] // U+9365 <cjk>
	`鍪`: [u8(0xEF), 0x5D] // U+936A <cjk>
	`鍰`: [u8(0xEF), 0x5E] // U+9370 <cjk>
	`鎛`: [u8(0xEF), 0x5F] // U+939B <cjk>
	`鎣`: [u8(0xEF), 0x60] // U+93A3 <cjk>
	`鎺`: [u8(0xEF), 0x61] // U+93BA <cjk>
	`鏆`: [u8(0xEF), 0x62] // U+93C6 <cjk>
	`鏞`: [u8(0xEF), 0x63] // U+93DE <cjk>
	`鏟`: [u8(0xEF), 0x64] // U+93DF <cjk>
	`鐄`: [u8(0xEF), 0x65] // U+9404 <cjk>
	`鏽`: [u8(0xEF), 0x66] // U+93FD <cjk>
	`鐳`: [u8(0xEF), 0x67] // U+9433 <cjk>
	`鑊`: [u8(0xEF), 0x68] // U+944A <cjk>
	`鑣`: [u8(0xEF), 0x69] // U+9463 <cjk>
	`鑫`: [u8(0xEF), 0x6A] // U+946B <cjk>
	`鑱`: [u8(0xEF), 0x6B] // U+9471 <cjk>
	`鑲`: [u8(0xEF), 0x6C] // U+9472 <cjk>
	`閎`: [u8(0xEF), 0x6D] // U+958E <cjk>
	`閟`: [u8(0xEF), 0x6E] // U+959F <cjk>
	`閦`: [u8(0xEF), 0x6F] // U+95A6 <cjk>
	`閩`: [u8(0xEF), 0x70] // U+95A9 <cjk>
	`閬`: [u8(0xEF), 0x71] // U+95AC <cjk>
	`閶`: [u8(0xEF), 0x72] // U+95B6 <cjk>
	`閽`: [u8(0xEF), 0x73] // U+95BD <cjk>
	`闋`: [u8(0xEF), 0x74] // U+95CB <cjk>
	`闐`: [u8(0xEF), 0x75] // U+95D0 <cjk>
	`闓`: [u8(0xEF), 0x76] // U+95D3 <cjk>
	`䦰`: [u8(0xEF), 0x77] // U+49B0 <cjk>
	`闚`: [u8(0xEF), 0x78] // U+95DA <cjk>
	`闞`: [u8(0xEF), 0x79] // U+95DE <cjk>
	`陘`: [u8(0xEF), 0x7A] // U+9658 <cjk>
	`隄`: [u8(0xEF), 0x7B] // U+9684 <cjk>
	`隆`: [u8(0xEF), 0x7C] // U+F9DC CJK COMPATIBILITY IDEOGRAPH-F9DC
	`隝`: [u8(0xEF), 0x7D] // U+969D <cjk>
	`隤`: [u8(0xEF), 0x7E] // U+96A4 <cjk>
	`隥`: [u8(0xEF), 0x80] // U+96A5 <cjk>
	`雒`: [u8(0xEF), 0x81] // U+96D2 <cjk>
	`雞`: [u8(0xEF), 0x82] // U+96DE <cjk>
	`難`: [u8(0xEF), 0x83] // U+FA68 CJK COMPATIBILITY IDEOGRAPH-FA68
	`雩`: [u8(0xEF), 0x84] // U+96E9 <cjk>
	`雯`: [u8(0xEF), 0x85] // U+96EF <cjk>
	`霳`: [u8(0xEF), 0x86] // U+9733 <cjk>
	`霻`: [u8(0xEF), 0x87] // U+973B <cjk>
	`靍`: [u8(0xEF), 0x88] // U+974D <cjk>
	`靎`: [u8(0xEF), 0x89] // U+974E <cjk>
	`靏`: [u8(0xEF), 0x8A] // U+974F <cjk>
	`靚`: [u8(0xEF), 0x8B] // U+975A <cjk>
	`靮`: [u8(0xEF), 0x8C] // U+976E <cjk>
	`靳`: [u8(0xEF), 0x8D] // U+9773 <cjk>
	`鞕`: [u8(0xEF), 0x8E] // U+9795 <cjk>
	`鞮`: [u8(0xEF), 0x8F] // U+97AE <cjk>
	`鞺`: [u8(0xEF), 0x90] // U+97BA <cjk>
	`韁`: [u8(0xEF), 0x91] // U+97C1 <cjk>
	`韉`: [u8(0xEF), 0x92] // U+97C9 <cjk>
	`韞`: [u8(0xEF), 0x93] // U+97DE <cjk>
	`韛`: [u8(0xEF), 0x94] // U+97DB <cjk>
	`韴`: [u8(0xEF), 0x95] // U+97F4 <cjk>
	`響`: [u8(0xEF), 0x96] // U+FA69 CJK COMPATIBILITY IDEOGRAPH-FA69
	`頊`: [u8(0xEF), 0x97] // U+980A <cjk>
	`頞`: [u8(0xEF), 0x98] // U+981E <cjk>
	`頫`: [u8(0xEF), 0x99] // U+982B <cjk>
	`頰`: [u8(0xEF), 0x9A] // U+9830 <cjk>
	`頻`: [u8(0xEF), 0x9B] // U+FA6A CJK COMPATIBILITY IDEOGRAPH-FA6A
	`顒`: [u8(0xEF), 0x9C] // U+9852 <cjk>
	`顓`: [u8(0xEF), 0x9D] // U+9853 <cjk>
	`顖`: [u8(0xEF), 0x9E] // U+9856 <cjk>
	`顗`: [u8(0xEF), 0x9F] // U+9857 <cjk>
	`顙`: [u8(0xEF), 0xA0] // U+9859 <cjk>
	`顚`: [u8(0xEF), 0xA1] // U+985A <cjk>
	`類`: [u8(0xEF), 0xA2] // U+F9D0 CJK COMPATIBILITY IDEOGRAPH-F9D0
	`顥`: [u8(0xEF), 0xA3] // U+9865 <cjk>
	`顬`: [u8(0xEF), 0xA4] // U+986C <cjk>
	`颺`: [u8(0xEF), 0xA5] // U+98BA <cjk>
	`飈`: [u8(0xEF), 0xA6] // U+98C8 <cjk>
	`飧`: [u8(0xEF), 0xA7] // U+98E7 <cjk>
	`饘`: [u8(0xEF), 0xA8] // U+9958 <cjk>
	`馞`: [u8(0xEF), 0xA9] // U+999E <cjk>
	`騂`: [u8(0xEF), 0xAA] // U+9A02 <cjk>
	`騃`: [u8(0xEF), 0xAB] // U+9A03 <cjk>
	`騤`: [u8(0xEF), 0xAC] // U+9A24 <cjk>
	`騭`: [u8(0xEF), 0xAD] // U+9A2D <cjk>
	`騮`: [u8(0xEF), 0xAE] // U+9A2E <cjk>
	`騸`: [u8(0xEF), 0xAF] // U+9A38 <cjk>
	`驊`: [u8(0xEF), 0xB0] // U+9A4A <cjk>
	`驎`: [u8(0xEF), 0xB1] // U+9A4E <cjk>
	`驒`: [u8(0xEF), 0xB2] // U+9A52 <cjk>
	`骶`: [u8(0xEF), 0xB3] // U+9AB6 <cjk>
	`髁`: [u8(0xEF), 0xB4] // U+9AC1 <cjk>
	`髃`: [u8(0xEF), 0xB5] // U+9AC3 <cjk>
	`髎`: [u8(0xEF), 0xB6] // U+9ACE <cjk>
	`髖`: [u8(0xEF), 0xB7] // U+9AD6 <cjk>
	`髹`: [u8(0xEF), 0xB8] // U+9AF9 <cjk>
	`鬂`: [u8(0xEF), 0xB9] // U+9B02 <cjk>
	`鬈`: [u8(0xEF), 0xBA] // U+9B08 <cjk>
	`鬠`: [u8(0xEF), 0xBB] // U+9B20 <cjk>
	`䰗`: [u8(0xEF), 0xBC] // U+4C17 <cjk>
	`鬭`: [u8(0xEF), 0xBD] // U+9B2D <cjk>
	`魞`: [u8(0xEF), 0xBE] // U+9B5E <cjk>
	`魹`: [u8(0xEF), 0xBF] // U+9B79 <cjk>
	`魦`: [u8(0xEF), 0xC0] // U+9B66 <cjk>
	`魲`: [u8(0xEF), 0xC1] // U+9B72 <cjk>
	`魵`: [u8(0xEF), 0xC2] // U+9B75 <cjk>
	`鮄`: [u8(0xEF), 0xC3] // U+9B84 <cjk>
	`鮊`: [u8(0xEF), 0xC4] // U+9B8A <cjk>
	`鮏`: [u8(0xEF), 0xC5] // U+9B8F <cjk>
	`鮞`: [u8(0xEF), 0xC6] // U+9B9E <cjk>
	`鮧`: [u8(0xEF), 0xC7] // U+9BA7 <cjk>
	`鯁`: [u8(0xEF), 0xC8] // U+9BC1 <cjk>
	`鯎`: [u8(0xEF), 0xC9] // U+9BCE <cjk>
	`鯥`: [u8(0xEF), 0xCA] // U+9BE5 <cjk>
	`鯸`: [u8(0xEF), 0xCB] // U+9BF8 <cjk>
	`鯽`: [u8(0xEF), 0xCC] // U+9BFD <cjk>
	`鰀`: [u8(0xEF), 0xCD] // U+9C00 <cjk>
	`鰣`: [u8(0xEF), 0xCE] // U+9C23 <cjk>
	`鱁`: [u8(0xEF), 0xCF] // U+9C41 <cjk>
	`鱏`: [u8(0xEF), 0xD0] // U+9C4F <cjk>
	`鱐`: [u8(0xEF), 0xD1] // U+9C50 <cjk>
	`鱓`: [u8(0xEF), 0xD2] // U+9C53 <cjk>
	`鱣`: [u8(0xEF), 0xD3] // U+9C63 <cjk>
	`鱥`: [u8(0xEF), 0xD4] // U+9C65 <cjk>
	`鱷`: [u8(0xEF), 0xD5] // U+9C77 <cjk>
	`鴝`: [u8(0xEF), 0xD6] // U+9D1D <cjk>
	`鴞`: [u8(0xEF), 0xD7] // U+9D1E <cjk>
	`鵃`: [u8(0xEF), 0xD8] // U+9D43 <cjk>
	`鵇`: [u8(0xEF), 0xD9] // U+9D47 <cjk>
	`鵒`: [u8(0xEF), 0xDA] // U+9D52 <cjk>
	`鵣`: [u8(0xEF), 0xDB] // U+9D63 <cjk>
	`鵰`: [u8(0xEF), 0xDC] // U+9D70 <cjk>
	`鵼`: [u8(0xEF), 0xDD] // U+9D7C <cjk>
	`鶊`: [u8(0xEF), 0xDE] // U+9D8A <cjk>
	`鶖`: [u8(0xEF), 0xDF] // U+9D96 <cjk>
	`鷀`: [u8(0xEF), 0xE0] // U+9DC0 <cjk>
	`鶬`: [u8(0xEF), 0xE1] // U+9DAC <cjk>
	`鶼`: [u8(0xEF), 0xE2] // U+9DBC <cjk>
	`鷗`: [u8(0xEF), 0xE3] // U+9DD7 <cjk>
	`𪆐`: [u8(0xEF), 0xE4] // U+2A190 <cjk>
	`鷧`: [u8(0xEF), 0xE5] // U+9DE7 <cjk>
	`鸇`: [u8(0xEF), 0xE6] // U+9E07 <cjk>
	`鸕`: [u8(0xEF), 0xE7] // U+9E15 <cjk>
	`鹼`: [u8(0xEF), 0xE8] // U+9E7C <cjk>
	`麞`: [u8(0xEF), 0xE9] // U+9E9E <cjk>
	`麤`: [u8(0xEF), 0xEA] // U+9EA4 <cjk>
	`麬`: [u8(0xEF), 0xEB] // U+9EAC <cjk>
	`麯`: [u8(0xEF), 0xEC] // U+9EAF <cjk>
	`麴`: [u8(0xEF), 0xED] // U+9EB4 <cjk>
	`麵`: [u8(0xEF), 0xEE] // U+9EB5 <cjk>
	`黃`: [u8(0xEF), 0xEF] // U+9EC3 <cjk>
	`黑`: [u8(0xEF), 0xF0] // U+9ED1 <cjk>
	`鼐`: [u8(0xEF), 0xF1] // U+9F10 <cjk>
	`鼹`: [u8(0xEF), 0xF2] // U+9F39 <cjk>
	`齗`: [u8(0xEF), 0xF3] // U+9F57 <cjk>
	`龐`: [u8(0xEF), 0xF4] // U+9F90 <cjk>
	`龔`: [u8(0xEF), 0xF5] // U+9F94 <cjk>
	`龗`: [u8(0xEF), 0xF6] // U+9F97 <cjk>
	`龢`: [u8(0xEF), 0xF7] // U+9FA2 <cjk>
	`姸`: [u8(0xEF), 0xF8] // U+59F8 <cjk>
	`屛`: [u8(0xEF), 0xF9] // U+5C5B <cjk>
	`幷`: [u8(0xEF), 0xFA] // U+5E77 <cjk>
	`瘦`: [u8(0xEF), 0xFB] // U+7626 <cjk>
	`繫`: [u8(0xEF), 0xFC] // U+7E6B <cjk>
	`𠂉`: [u8(0xF0), 0x40] // U+20089 <cjk>
	`丂`: [u8(0xF0), 0x41] // U+4E02 <cjk>
	`丏`: [u8(0xF0), 0x42] // U+4E0F <cjk>
	`丒`: [u8(0xF0), 0x43] // U+4E12 <cjk>
	`丩`: [u8(0xF0), 0x44] // U+4E29 <cjk>
	`丫`: [u8(0xF0), 0x45] // U+4E2B <cjk>
	`丮`: [u8(0xF0), 0x46] // U+4E2E <cjk>
	`乀`: [u8(0xF0), 0x47] // U+4E40 <cjk>
	`乇`: [u8(0xF0), 0x48] // U+4E47 <cjk>
	`么`: [u8(0xF0), 0x49] // U+4E48 <cjk>
	`𠂢`: [u8(0xF0), 0x4A] // U+200A2 <cjk>
	`乑`: [u8(0xF0), 0x4B] // U+4E51 <cjk>
	`㐆`: [u8(0xF0), 0x4C] // U+3406 <cjk>
	`𠂤`: [u8(0xF0), 0x4D] // U+200A4 <cjk>
	`乚`: [u8(0xF0), 0x4E] // U+4E5A <cjk>
	`乩`: [u8(0xF0), 0x4F] // U+4E69 <cjk>
	`亝`: [u8(0xF0), 0x50] // U+4E9D <cjk>
	`㐬`: [u8(0xF0), 0x51] // U+342C <cjk>
	`㐮`: [u8(0xF0), 0x52] // U+342E <cjk>
	`亹`: [u8(0xF0), 0x53] // U+4EB9 <cjk>
	`亻`: [u8(0xF0), 0x54] // U+4EBB <cjk>
	`𠆢`: [u8(0xF0), 0x55] // U+201A2 <cjk>
	`亼`: [u8(0xF0), 0x56] // U+4EBC <cjk>
	`仃`: [u8(0xF0), 0x57] // U+4EC3 <cjk>
	`仈`: [u8(0xF0), 0x58] // U+4EC8 <cjk>
	`仐`: [u8(0xF0), 0x59] // U+4ED0 <cjk>
	`仫`: [u8(0xF0), 0x5A] // U+4EEB <cjk>
	`仚`: [u8(0xF0), 0x5B] // U+4EDA <cjk>
	`仱`: [u8(0xF0), 0x5C] // U+4EF1 <cjk>
	`仵`: [u8(0xF0), 0x5D] // U+4EF5 <cjk>
	`伀`: [u8(0xF0), 0x5E] // U+4F00 <cjk>
	`伖`: [u8(0xF0), 0x5F] // U+4F16 <cjk>
	`佤`: [u8(0xF0), 0x60] // U+4F64 <cjk>
	`伷`: [u8(0xF0), 0x61] // U+4F37 <cjk>
	`伾`: [u8(0xF0), 0x62] // U+4F3E <cjk>
	`佔`: [u8(0xF0), 0x63] // U+4F54 <cjk>
	`佘`: [u8(0xF0), 0x64] // U+4F58 <cjk>
	`𠈓`: [u8(0xF0), 0x65] // U+20213 <cjk>
	`佷`: [u8(0xF0), 0x66] // U+4F77 <cjk>
	`佸`: [u8(0xF0), 0x67] // U+4F78 <cjk>
	`佺`: [u8(0xF0), 0x68] // U+4F7A <cjk>
	`佽`: [u8(0xF0), 0x69] // U+4F7D <cjk>
	`侂`: [u8(0xF0), 0x6A] // U+4F82 <cjk>
	`侅`: [u8(0xF0), 0x6B] // U+4F85 <cjk>
	`侒`: [u8(0xF0), 0x6C] // U+4F92 <cjk>
	`侚`: [u8(0xF0), 0x6D] // U+4F9A <cjk>
	`俦`: [u8(0xF0), 0x6E] // U+4FE6 <cjk>
	`侲`: [u8(0xF0), 0x6F] // U+4FB2 <cjk>
	`侾`: [u8(0xF0), 0x70] // U+4FBE <cjk>
	`俅`: [u8(0xF0), 0x71] // U+4FC5 <cjk>
	`俋`: [u8(0xF0), 0x72] // U+4FCB <cjk>
	`俏`: [u8(0xF0), 0x73] // U+4FCF <cjk>
	`俒`: [u8(0xF0), 0x74] // U+4FD2 <cjk>
	`㑪`: [u8(0xF0), 0x75] // U+346A <cjk>
	`俲`: [u8(0xF0), 0x76] // U+4FF2 <cjk>
	`倀`: [u8(0xF0), 0x77] // U+5000 <cjk>
	`倐`: [u8(0xF0), 0x78] // U+5010 <cjk>
	`倓`: [u8(0xF0), 0x79] // U+5013 <cjk>
	`倜`: [u8(0xF0), 0x7A] // U+501C <cjk>
	`倞`: [u8(0xF0), 0x7B] // U+501E <cjk>
	`倢`: [u8(0xF0), 0x7C] // U+5022 <cjk>
	`㑨`: [u8(0xF0), 0x7D] // U+3468 <cjk>
	`偂`: [u8(0xF0), 0x7E] // U+5042 <cjk>
	`偆`: [u8(0xF0), 0x80] // U+5046 <cjk>
	`偎`: [u8(0xF0), 0x81] // U+504E <cjk>
	`偓`: [u8(0xF0), 0x82] // U+5053 <cjk>
	`偗`: [u8(0xF0), 0x83] // U+5057 <cjk>
	`偣`: [u8(0xF0), 0x84] // U+5063 <cjk>
	`偦`: [u8(0xF0), 0x85] // U+5066 <cjk>
	`偪`: [u8(0xF0), 0x86] // U+506A <cjk>
	`偰`: [u8(0xF0), 0x87] // U+5070 <cjk>
	`傣`: [u8(0xF0), 0x88] // U+50A3 <cjk>
	`傈`: [u8(0xF0), 0x89] // U+5088 <cjk>
	`傒`: [u8(0xF0), 0x8A] // U+5092 <cjk>
	`傓`: [u8(0xF0), 0x8B] // U+5093 <cjk>
	`傕`: [u8(0xF0), 0x8C] // U+5095 <cjk>
	`傖`: [u8(0xF0), 0x8D] // U+5096 <cjk>
	`傜`: [u8(0xF0), 0x8E] // U+509C <cjk>
	`傪`: [u8(0xF0), 0x8F] // U+50AA <cjk>
	`𠌫`: [u8(0xF0), 0x90] // U+2032B <cjk>
	`傱`: [u8(0xF0), 0x91] // U+50B1 <cjk>
	`傺`: [u8(0xF0), 0x92] // U+50BA <cjk>
	`傻`: [u8(0xF0), 0x93] // U+50BB <cjk>
	`僄`: [u8(0xF0), 0x94] // U+50C4 <cjk>
	`僇`: [u8(0xF0), 0x95] // U+50C7 <cjk>
	`僳`: [u8(0xF0), 0x96] // U+50F3 <cjk>
	`𠎁`: [u8(0xF0), 0x97] // U+20381 <cjk>
	`僎`: [u8(0xF0), 0x98] // U+50CE <cjk>
	`𠍱`: [u8(0xF0), 0x99] // U+20371 <cjk>
	`僔`: [u8(0xF0), 0x9A] // U+50D4 <cjk>
	`僙`: [u8(0xF0), 0x9B] // U+50D9 <cjk>
	`僡`: [u8(0xF0), 0x9C] // U+50E1 <cjk>
	`僩`: [u8(0xF0), 0x9D] // U+50E9 <cjk>
	`㒒`: [u8(0xF0), 0x9E] // U+3492 <cjk>
	`宖`: [u8(0xF0), 0x9F] // U+5B96 <cjk>
	`宬`: [u8(0xF0), 0xA0] // U+5BAC <cjk>
	`㝡`: [u8(0xF0), 0xA1] // U+3761 <cjk>
	`寀`: [u8(0xF0), 0xA2] // U+5BC0 <cjk>
	`㝢`: [u8(0xF0), 0xA3] // U+3762 <cjk>
	`寎`: [u8(0xF0), 0xA4] // U+5BCE <cjk>
	`寖`: [u8(0xF0), 0xA5] // U+5BD6 <cjk>
	`㝬`: [u8(0xF0), 0xA6] // U+376C <cjk>
	`㝫`: [u8(0xF0), 0xA7] // U+376B <cjk>
	`寱`: [u8(0xF0), 0xA8] // U+5BF1 <cjk>
	`寽`: [u8(0xF0), 0xA9] // U+5BFD <cjk>
	`㝵`: [u8(0xF0), 0xAA] // U+3775 <cjk>
	`尃`: [u8(0xF0), 0xAB] // U+5C03 <cjk>
	`尩`: [u8(0xF0), 0xAC] // U+5C29 <cjk>
	`尰`: [u8(0xF0), 0xAD] // U+5C30 <cjk>
	`𡱖`: [u8(0xF0), 0xAE] // U+21C56 <cjk>
	`屟`: [u8(0xF0), 0xAF] // U+5C5F <cjk>
	`屣`: [u8(0xF0), 0xB0] // U+5C63 <cjk>
	`屧`: [u8(0xF0), 0xB1] // U+5C67 <cjk>
	`屨`: [u8(0xF0), 0xB2] // U+5C68 <cjk>
	`屩`: [u8(0xF0), 0xB3] // U+5C69 <cjk>
	`屰`: [u8(0xF0), 0xB4] // U+5C70 <cjk>
	`𡴭`: [u8(0xF0), 0xB5] // U+21D2D <cjk>
	`𡵅`: [u8(0xF0), 0xB6] // U+21D45 <cjk>
	`屼`: [u8(0xF0), 0xB7] // U+5C7C <cjk>
	`𡵸`: [u8(0xF0), 0xB8] // U+21D78 <cjk>
	`𡵢`: [u8(0xF0), 0xB9] // U+21D62 <cjk>
	`岈`: [u8(0xF0), 0xBA] // U+5C88 <cjk>
	`岊`: [u8(0xF0), 0xBB] // U+5C8A <cjk>
	`㟁`: [u8(0xF0), 0xBC] // U+37C1 <cjk>
	`𡶡`: [u8(0xF0), 0xBD] // U+21DA1 <cjk>
	`𡶜`: [u8(0xF0), 0xBE] // U+21D9C <cjk>
	`岠`: [u8(0xF0), 0xBF] // U+5CA0 <cjk>
	`岢`: [u8(0xF0), 0xC0] // U+5CA2 <cjk>
	`岦`: [u8(0xF0), 0xC1] // U+5CA6 <cjk>
	`岧`: [u8(0xF0), 0xC2] // U+5CA7 <cjk>
	`𡶒`: [u8(0xF0), 0xC3] // U+21D92 <cjk>
	`岭`: [u8(0xF0), 0xC4] // U+5CAD <cjk>
	`岵`: [u8(0xF0), 0xC5] // U+5CB5 <cjk>
	`𡶷`: [u8(0xF0), 0xC6] // U+21DB7 <cjk>
	`峉`: [u8(0xF0), 0xC7] // U+5CC9 <cjk>
	`𡷠`: [u8(0xF0), 0xC8] // U+21DE0 <cjk>
	`𡸳`: [u8(0xF0), 0xC9] // U+21E33 <cjk>
	`崆`: [u8(0xF0), 0xCA] // U+5D06 <cjk>
	`崐`: [u8(0xF0), 0xCB] // U+5D10 <cjk>
	`崫`: [u8(0xF0), 0xCC] // U+5D2B <cjk>
	`崝`: [u8(0xF0), 0xCD] // U+5D1D <cjk>
	`崠`: [u8(0xF0), 0xCE] // U+5D20 <cjk>
	`崤`: [u8(0xF0), 0xCF] // U+5D24 <cjk>
	`崦`: [u8(0xF0), 0xD0] // U+5D26 <cjk>
	`崱`: [u8(0xF0), 0xD1] // U+5D31 <cjk>
	`崹`: [u8(0xF0), 0xD2] // U+5D39 <cjk>
	`嵂`: [u8(0xF0), 0xD3] // U+5D42 <cjk>
	`㟨`: [u8(0xF0), 0xD4] // U+37E8 <cjk>
	`嵡`: [u8(0xF0), 0xD5] // U+5D61 <cjk>
	`嵪`: [u8(0xF0), 0xD6] // U+5D6A <cjk>
	`㟴`: [u8(0xF0), 0xD7] // U+37F4 <cjk>
	`嵰`: [u8(0xF0), 0xD8] // U+5D70 <cjk>
	`𡼞`: [u8(0xF0), 0xD9] // U+21F1E <cjk>
	`㟽`: [u8(0xF0), 0xDA] // U+37FD <cjk>
	`嶈`: [u8(0xF0), 0xDB] // U+5D88 <cjk>
	`㠀`: [u8(0xF0), 0xDC] // U+3800 <cjk>
	`嶒`: [u8(0xF0), 0xDD] // U+5D92 <cjk>
	`嶔`: [u8(0xF0), 0xDE] // U+5D94 <cjk>
	`嶗`: [u8(0xF0), 0xDF] // U+5D97 <cjk>
	`嶙`: [u8(0xF0), 0xE0] // U+5D99 <cjk>
	`嶰`: [u8(0xF0), 0xE1] // U+5DB0 <cjk>
	`嶲`: [u8(0xF0), 0xE2] // U+5DB2 <cjk>
	`嶴`: [u8(0xF0), 0xE3] // U+5DB4 <cjk>
	`𡽶`: [u8(0xF0), 0xE4] // U+21F76 <cjk>
	`嶹`: [u8(0xF0), 0xE5] // U+5DB9 <cjk>
	`巑`: [u8(0xF0), 0xE6] // U+5DD1 <cjk>
	`巗`: [u8(0xF0), 0xE7] // U+5DD7 <cjk>
	`巘`: [u8(0xF0), 0xE8] // U+5DD8 <cjk>
	`巠`: [u8(0xF0), 0xE9] // U+5DE0 <cjk>
	`𡿺`: [u8(0xF0), 0xEA] // U+21FFA <cjk>
	`巤`: [u8(0xF0), 0xEB] // U+5DE4 <cjk>
	`巩`: [u8(0xF0), 0xEC] // U+5DE9 <cjk>
	`㠯`: [u8(0xF0), 0xED] // U+382F <cjk>
	`帀`: [u8(0xF0), 0xEE] // U+5E00 <cjk>
	`㠶`: [u8(0xF0), 0xEF] // U+3836 <cjk>
	`帒`: [u8(0xF0), 0xF0] // U+5E12 <cjk>
	`帕`: [u8(0xF0), 0xF1] // U+5E15 <cjk>
	`㡀`: [u8(0xF0), 0xF2] // U+3840 <cjk>
	`帟`: [u8(0xF0), 0xF3] // U+5E1F <cjk>
	`帮`: [u8(0xF0), 0xF4] // U+5E2E <cjk>
	`帾`: [u8(0xF0), 0xF5] // U+5E3E <cjk>
	`幉`: [u8(0xF0), 0xF6] // U+5E49 <cjk>
	`㡜`: [u8(0xF0), 0xF7] // U+385C <cjk>
	`幖`: [u8(0xF0), 0xF8] // U+5E56 <cjk>
	`㡡`: [u8(0xF0), 0xF9] // U+3861 <cjk>
	`幫`: [u8(0xF0), 0xFA] // U+5E6B <cjk>
	`幬`: [u8(0xF0), 0xFB] // U+5E6C <cjk>
	`幭`: [u8(0xF0), 0xFC] // U+5E6D <cjk>
	`儈`: [u8(0xF1), 0x40] // U+5108 <cjk>
	`𠏹`: [u8(0xF1), 0x41] // U+203F9 <cjk>
	`儗`: [u8(0xF1), 0x42] // U+5117 <cjk>
	`儛`: [u8(0xF1), 0x43] // U+511B <cjk>
	`𠑊`: [u8(0xF1), 0x44] // U+2044A <cjk>
	`兠`: [u8(0xF1), 0x45] // U+5160 <cjk>
	`𠔉`: [u8(0xF1), 0x46] // U+20509 <cjk>
	`关`: [u8(0xF1), 0x47] // U+5173 <cjk>
	`冃`: [u8(0xF1), 0x48] // U+5183 <cjk>
	`冋`: [u8(0xF1), 0x49] // U+518B <cjk>
	`㒼`: [u8(0xF1), 0x4A] // U+34BC <cjk>
	`冘`: [u8(0xF1), 0x4B] // U+5198 <cjk>
	`冣`: [u8(0xF1), 0x4C] // U+51A3 <cjk>
	`冭`: [u8(0xF1), 0x4D] // U+51AD <cjk>
	`㓇`: [u8(0xF1), 0x4E] // U+34C7 <cjk>
	`冼`: [u8(0xF1), 0x4F] // U+51BC <cjk>
	`𠗖`: [u8(0xF1), 0x50] // U+205D6 <cjk>
	`𠘨`: [u8(0xF1), 0x51] // U+20628 <cjk>
	`凳`: [u8(0xF1), 0x52] // U+51F3 <cjk>
	`凴`: [u8(0xF1), 0x53] // U+51F4 <cjk>
	`刂`: [u8(0xF1), 0x54] // U+5202 <cjk>
	`划`: [u8(0xF1), 0x55] // U+5212 <cjk>
	`刖`: [u8(0xF1), 0x56] // U+5216 <cjk>
	`𠝏`: [u8(0xF1), 0x57] // U+2074F <cjk>
	`剕`: [u8(0xF1), 0x58] // U+5255 <cjk>
	`剜`: [u8(0xF1), 0x59] // U+525C <cjk>
	`剬`: [u8(0xF1), 0x5A] // U+526C <cjk>
	`剷`: [u8(0xF1), 0x5B] // U+5277 <cjk>
	`劄`: [u8(0xF1), 0x5C] // U+5284 <cjk>
	`劂`: [u8(0xF1), 0x5D] // U+5282 <cjk>
	`𠠇`: [u8(0xF1), 0x5E] // U+20807 <cjk>
	`劘`: [u8(0xF1), 0x5F] // U+5298 <cjk>
	`𠠺`: [u8(0xF1), 0x60] // U+2083A <cjk>
	`劤`: [u8(0xF1), 0x61] // U+52A4 <cjk>
	`劦`: [u8(0xF1), 0x62] // U+52A6 <cjk>
	`劯`: [u8(0xF1), 0x63] // U+52AF <cjk>
	`劺`: [u8(0xF1), 0x64] // U+52BA <cjk>
	`劻`: [u8(0xF1), 0x65] // U+52BB <cjk>
	`勊`: [u8(0xF1), 0x66] // U+52CA <cjk>
	`㔟`: [u8(0xF1), 0x67] // U+351F <cjk>
	`勑`: [u8(0xF1), 0x68] // U+52D1 <cjk>
	`𠢹`: [u8(0xF1), 0x69] // U+208B9 <cjk>
	`勷`: [u8(0xF1), 0x6A] // U+52F7 <cjk>
	`匊`: [u8(0xF1), 0x6B] // U+530A <cjk>
	`匋`: [u8(0xF1), 0x6C] // U+530B <cjk>
	`匤`: [u8(0xF1), 0x6D] // U+5324 <cjk>
	`匵`: [u8(0xF1), 0x6E] // U+5335 <cjk>
	`匾`: [u8(0xF1), 0x6F] // U+533E <cjk>
	`卂`: [u8(0xF1), 0x70] // U+5342 <cjk>
	`𠥼`: [u8(0xF1), 0x71] // U+2097C <cjk>
	`𠦝`: [u8(0xF1), 0x72] // U+2099D <cjk>
	`卧`: [u8(0xF1), 0x73] // U+5367 <cjk>
	`卬`: [u8(0xF1), 0x74] // U+536C <cjk>
	`卺`: [u8(0xF1), 0x75] // U+537A <cjk>
	`厤`: [u8(0xF1), 0x76] // U+53A4 <cjk>
	`厴`: [u8(0xF1), 0x77] // U+53B4 <cjk>
	`𠫓`: [u8(0xF1), 0x78] // U+20AD3 <cjk>
	`厷`: [u8(0xF1), 0x79] // U+53B7 <cjk>
	`叀`: [u8(0xF1), 0x7A] // U+53C0 <cjk>
	`𠬝`: [u8(0xF1), 0x7B] // U+20B1D <cjk>
	`㕝`: [u8(0xF1), 0x7C] // U+355D <cjk>
	`㕞`: [u8(0xF1), 0x7D] // U+355E <cjk>
	`叕`: [u8(0xF1), 0x7E] // U+53D5 <cjk>
	`叚`: [u8(0xF1), 0x80] // U+53DA <cjk>
	`㕣`: [u8(0xF1), 0x81] // U+3563 <cjk>
	`叴`: [u8(0xF1), 0x82] // U+53F4 <cjk>
	`叵`: [u8(0xF1), 0x83] // U+53F5 <cjk>
	`呕`: [u8(0xF1), 0x84] // U+5455 <cjk>
	`吤`: [u8(0xF1), 0x85] // U+5424 <cjk>
	`吨`: [u8(0xF1), 0x86] // U+5428 <cjk>
	`㕮`: [u8(0xF1), 0x87] // U+356E <cjk>
	`呃`: [u8(0xF1), 0x88] // U+5443 <cjk>
	`呢`: [u8(0xF1), 0x89] // U+5462 <cjk>
	`呦`: [u8(0xF1), 0x8A] // U+5466 <cjk>
	`呬`: [u8(0xF1), 0x8B] // U+546C <cjk>
	`咊`: [u8(0xF1), 0x8C] // U+548A <cjk>
	`咍`: [u8(0xF1), 0x8D] // U+548D <cjk>
	`咕`: [u8(0xF1), 0x8E] // U+5495 <cjk>
	`咠`: [u8(0xF1), 0x8F] // U+54A0 <cjk>
	`咦`: [u8(0xF1), 0x90] // U+54A6 <cjk>
	`咭`: [u8(0xF1), 0x91] // U+54AD <cjk>
	`咮`: [u8(0xF1), 0x92] // U+54AE <cjk>
	`咷`: [u8(0xF1), 0x93] // U+54B7 <cjk>
	`咺`: [u8(0xF1), 0x94] // U+54BA <cjk>
	`咿`: [u8(0xF1), 0x95] // U+54BF <cjk>
	`哃`: [u8(0xF1), 0x96] // U+54C3 <cjk>
	`𠵅`: [u8(0xF1), 0x97] // U+20D45 <cjk>
	`哬`: [u8(0xF1), 0x98] // U+54EC <cjk>
	`哯`: [u8(0xF1), 0x99] // U+54EF <cjk>
	`哱`: [u8(0xF1), 0x9A] // U+54F1 <cjk>
	`哳`: [u8(0xF1), 0x9B] // U+54F3 <cjk>
	`唀`: [u8(0xF1), 0x9C] // U+5500 <cjk>
	`唁`: [u8(0xF1), 0x9D] // U+5501 <cjk>
	`唉`: [u8(0xF1), 0x9E] // U+5509 <cjk>
	`唼`: [u8(0xF1), 0x9F] // U+553C <cjk>
	`啁`: [u8(0xF1), 0xA0] // U+5541 <cjk>
	`㖦`: [u8(0xF1), 0xA1] // U+35A6 <cjk>
	`啇`: [u8(0xF1), 0xA2] // U+5547 <cjk>
	`啊`: [u8(0xF1), 0xA3] // U+554A <cjk>
	`㖨`: [u8(0xF1), 0xA4] // U+35A8 <cjk>
	`啠`: [u8(0xF1), 0xA5] // U+5560 <cjk>
	`啡`: [u8(0xF1), 0xA6] // U+5561 <cjk>
	`啤`: [u8(0xF1), 0xA7] // U+5564 <cjk>
	`𠷡`: [u8(0xF1), 0xA8] // U+20DE1 <cjk>
	`啽`: [u8(0xF1), 0xA9] // U+557D <cjk>
	`喂`: [u8(0xF1), 0xAA] // U+5582 <cjk>
	`喈`: [u8(0xF1), 0xAB] // U+5588 <cjk>
	`喑`: [u8(0xF1), 0xAC] // U+5591 <cjk>
	`㗅`: [u8(0xF1), 0xAD] // U+35C5 <cjk>
	`嗒`: [u8(0xF1), 0xAE] // U+55D2 <cjk>
	`𠺕`: [u8(0xF1), 0xAF] // U+20E95 <cjk>
	`𠹭`: [u8(0xF1), 0xB0] // U+20E6D <cjk>
	`喿`: [u8(0xF1), 0xB1] // U+55BF <cjk>
	`嗉`: [u8(0xF1), 0xB2] // U+55C9 <cjk>
	`嗌`: [u8(0xF1), 0xB3] // U+55CC <cjk>
	`嗑`: [u8(0xF1), 0xB4] // U+55D1 <cjk>
	`嗝`: [u8(0xF1), 0xB5] // U+55DD <cjk>
	`㗚`: [u8(0xF1), 0xB6] // U+35DA <cjk>
	`嗢`: [u8(0xF1), 0xB7] // U+55E2 <cjk>
	`𠹤`: [u8(0xF1), 0xB8] // U+20E64 <cjk>
	`嗩`: [u8(0xF1), 0xB9] // U+55E9 <cjk>
	`嘨`: [u8(0xF1), 0xBA] // U+5628 <cjk>
	`𠽟`: [u8(0xF1), 0xBB] // U+20F5F <cjk>
	`嘇`: [u8(0xF1), 0xBC] // U+5607 <cjk>
	`嘐`: [u8(0xF1), 0xBD] // U+5610 <cjk>
	`嘰`: [u8(0xF1), 0xBE] // U+5630 <cjk>
	`嘷`: [u8(0xF1), 0xBF] // U+5637 <cjk>
	`㗴`: [u8(0xF1), 0xC0] // U+35F4 <cjk>
	`嘽`: [u8(0xF1), 0xC1] // U+563D <cjk>
	`嘿`: [u8(0xF1), 0xC2] // U+563F <cjk>
	`噀`: [u8(0xF1), 0xC3] // U+5640 <cjk>
	`噇`: [u8(0xF1), 0xC4] // U+5647 <cjk>
	`噞`: [u8(0xF1), 0xC5] // U+565E <cjk>
	`噠`: [u8(0xF1), 0xC6] // U+5660 <cjk>
	`噭`: [u8(0xF1), 0xC7] // U+566D <cjk>
	`㘅`: [u8(0xF1), 0xC8] // U+3605 <cjk>
	`嚈`: [u8(0xF1), 0xC9] // U+5688 <cjk>
	`嚌`: [u8(0xF1), 0xCA] // U+568C <cjk>
	`嚕`: [u8(0xF1), 0xCB] // U+5695 <cjk>
	`嚚`: [u8(0xF1), 0xCC] // U+569A <cjk>
	`嚝`: [u8(0xF1), 0xCD] // U+569D <cjk>
	`嚨`: [u8(0xF1), 0xCE] // U+56A8 <cjk>
	`嚭`: [u8(0xF1), 0xCF] // U+56AD <cjk>
	`嚲`: [u8(0xF1), 0xD0] // U+56B2 <cjk>
	`囅`: [u8(0xF1), 0xD1] // U+56C5 <cjk>
	`囍`: [u8(0xF1), 0xD2] // U+56CD <cjk>
	`囟`: [u8(0xF1), 0xD3] // U+56DF <cjk>
	`囨`: [u8(0xF1), 0xD4] // U+56E8 <cjk>
	`囶`: [u8(0xF1), 0xD5] // U+56F6 <cjk>
	`囷`: [u8(0xF1), 0xD6] // U+56F7 <cjk>
	`𡈁`: [u8(0xF1), 0xD7] // U+21201 <cjk>
	`圕`: [u8(0xF1), 0xD8] // U+5715 <cjk>
	`圣`: [u8(0xF1), 0xD9] // U+5723 <cjk>
	`𡉕`: [u8(0xF1), 0xDA] // U+21255 <cjk>
	`圩`: [u8(0xF1), 0xDB] // U+5729 <cjk>
	`𡉻`: [u8(0xF1), 0xDC] // U+2127B <cjk>
	`坅`: [u8(0xF1), 0xDD] // U+5745 <cjk>
	`坆`: [u8(0xF1), 0xDE] // U+5746 <cjk>
	`坌`: [u8(0xF1), 0xDF] // U+574C <cjk>
	`坍`: [u8(0xF1), 0xE0] // U+574D <cjk>
	`𡉴`: [u8(0xF1), 0xE1] // U+21274 <cjk>
	`坨`: [u8(0xF1), 0xE2] // U+5768 <cjk>
	`坯`: [u8(0xF1), 0xE3] // U+576F <cjk>
	`坳`: [u8(0xF1), 0xE4] // U+5773 <cjk>
	`坴`: [u8(0xF1), 0xE5] // U+5774 <cjk>
	`坵`: [u8(0xF1), 0xE6] // U+5775 <cjk>
	`坻`: [u8(0xF1), 0xE7] // U+577B <cjk>
	`𡋤`: [u8(0xF1), 0xE8] // U+212E4 <cjk>
	`𡋗`: [u8(0xF1), 0xE9] // U+212D7 <cjk>
	`垬`: [u8(0xF1), 0xEA] // U+57AC <cjk>
	`垚`: [u8(0xF1), 0xEB] // U+579A <cjk>
	`垝`: [u8(0xF1), 0xEC] // U+579D <cjk>
	`垞`: [u8(0xF1), 0xED] // U+579E <cjk>
	`垨`: [u8(0xF1), 0xEE] // U+57A8 <cjk>
	`埗`: [u8(0xF1), 0xEF] // U+57D7 <cjk>
	`𡋽`: [u8(0xF1), 0xF0] // U+212FD <cjk>
	`埌`: [u8(0xF1), 0xF1] // U+57CC <cjk>
	`𡌶`: [u8(0xF1), 0xF2] // U+21336 <cjk>
	`𡍄`: [u8(0xF1), 0xF3] // U+21344 <cjk>
	`埞`: [u8(0xF1), 0xF4] // U+57DE <cjk>
	`埦`: [u8(0xF1), 0xF5] // U+57E6 <cjk>
	`埰`: [u8(0xF1), 0xF6] // U+57F0 <cjk>
	`㙊`: [u8(0xF1), 0xF7] // U+364A <cjk>
	`埸`: [u8(0xF1), 0xF8] // U+57F8 <cjk>
	`埻`: [u8(0xF1), 0xF9] // U+57FB <cjk>
	`埽`: [u8(0xF1), 0xFA] // U+57FD <cjk>
	`堄`: [u8(0xF1), 0xFB] // U+5804 <cjk>
	`堞`: [u8(0xF1), 0xFC] // U+581E <cjk>
	`堠`: [u8(0xF2), 0x40] // U+5820 <cjk>
	`堧`: [u8(0xF2), 0x41] // U+5827 <cjk>
	`堲`: [u8(0xF2), 0x42] // U+5832 <cjk>
	`堹`: [u8(0xF2), 0x43] // U+5839 <cjk>
	`𡏄`: [u8(0xF2), 0x44] // U+213C4 <cjk>
	`塉`: [u8(0xF2), 0x45] // U+5849 <cjk>
	`塌`: [u8(0xF2), 0x46] // U+584C <cjk>
	`塧`: [u8(0xF2), 0x47] // U+5867 <cjk>
	`墊`: [u8(0xF2), 0x48] // U+588A <cjk>
	`墋`: [u8(0xF2), 0x49] // U+588B <cjk>
	`墍`: [u8(0xF2), 0x4A] // U+588D <cjk>
	`墏`: [u8(0xF2), 0x4B] // U+588F <cjk>
	`墐`: [u8(0xF2), 0x4C] // U+5890 <cjk>
	`墔`: [u8(0xF2), 0x4D] // U+5894 <cjk>
	`墝`: [u8(0xF2), 0x4E] // U+589D <cjk>
	`墪`: [u8(0xF2), 0x4F] // U+58AA <cjk>
	`墱`: [u8(0xF2), 0x50] // U+58B1 <cjk>
	`𡑭`: [u8(0xF2), 0x51] // U+2146D <cjk>
	`壃`: [u8(0xF2), 0x52] // U+58C3 <cjk>
	`壍`: [u8(0xF2), 0x53] // U+58CD <cjk>
	`壢`: [u8(0xF2), 0x54] // U+58E2 <cjk>
	`壳`: [u8(0xF2), 0x55] // U+58F3 <cjk>
	`壴`: [u8(0xF2), 0x56] // U+58F4 <cjk>
	`夅`: [u8(0xF2), 0x57] // U+5905 <cjk>
	`夆`: [u8(0xF2), 0x58] // U+5906 <cjk>
	`夋`: [u8(0xF2), 0x59] // U+590B <cjk>
	`复`: [u8(0xF2), 0x5A] // U+590D <cjk>
	`夔`: [u8(0xF2), 0x5B] // U+5914 <cjk>
	`夤`: [u8(0xF2), 0x5C] // U+5924 <cjk>
	`𡗗`: [u8(0xF2), 0x5D] // U+215D7 <cjk>
	`㚑`: [u8(0xF2), 0x5E] // U+3691 <cjk>
	`夽`: [u8(0xF2), 0x5F] // U+593D <cjk>
	`㚙`: [u8(0xF2), 0x60] // U+3699 <cjk>
	`奆`: [u8(0xF2), 0x61] // U+5946 <cjk>
	`㚖`: [u8(0xF2), 0x62] // U+3696 <cjk>
	`𦰩`: [u8(0xF2), 0x63] // U+26C29 <cjk>
	`奛`: [u8(0xF2), 0x64] // U+595B <cjk>
	`奟`: [u8(0xF2), 0x65] // U+595F <cjk>
	`𡙇`: [u8(0xF2), 0x66] // U+21647 <cjk>
	`奵`: [u8(0xF2), 0x67] // U+5975 <cjk>
	`奶`: [u8(0xF2), 0x68] // U+5976 <cjk>
	`奼`: [u8(0xF2), 0x69] // U+597C <cjk>
	`妟`: [u8(0xF2), 0x6A] // U+599F <cjk>
	`妮`: [u8(0xF2), 0x6B] // U+59AE <cjk>
	`妼`: [u8(0xF2), 0x6C] // U+59BC <cjk>
	`姈`: [u8(0xF2), 0x6D] // U+59C8 <cjk>
	`姍`: [u8(0xF2), 0x6E] // U+59CD <cjk>
	`姞`: [u8(0xF2), 0x6F] // U+59DE <cjk>
	`姣`: [u8(0xF2), 0x70] // U+59E3 <cjk>
	`姤`: [u8(0xF2), 0x71] // U+59E4 <cjk>
	`姧`: [u8(0xF2), 0x72] // U+59E7 <cjk>
	`姮`: [u8(0xF2), 0x73] // U+59EE <cjk>
	`𡜆`: [u8(0xF2), 0x74] // U+21706 <cjk>
	`𡝂`: [u8(0xF2), 0x75] // U+21742 <cjk>
	`㛏`: [u8(0xF2), 0x76] // U+36CF <cjk>
	`娌`: [u8(0xF2), 0x77] // U+5A0C <cjk>
	`娍`: [u8(0xF2), 0x78] // U+5A0D <cjk>
	`娗`: [u8(0xF2), 0x79] // U+5A17 <cjk>
	`娧`: [u8(0xF2), 0x7A] // U+5A27 <cjk>
	`娭`: [u8(0xF2), 0x7B] // U+5A2D <cjk>
	`婕`: [u8(0xF2), 0x7C] // U+5A55 <cjk>
	`婥`: [u8(0xF2), 0x7D] // U+5A65 <cjk>
	`婺`: [u8(0xF2), 0x7E] // U+5A7A <cjk>
	`媋`: [u8(0xF2), 0x80] // U+5A8B <cjk>
	`媜`: [u8(0xF2), 0x81] // U+5A9C <cjk>
	`媟`: [u8(0xF2), 0x82] // U+5A9F <cjk>
	`媠`: [u8(0xF2), 0x83] // U+5AA0 <cjk>
	`媢`: [u8(0xF2), 0x84] // U+5AA2 <cjk>
	`媱`: [u8(0xF2), 0x85] // U+5AB1 <cjk>
	`媳`: [u8(0xF2), 0x86] // U+5AB3 <cjk>
	`媵`: [u8(0xF2), 0x87] // U+5AB5 <cjk>
	`媺`: [u8(0xF2), 0x88] // U+5ABA <cjk>
	`媿`: [u8(0xF2), 0x89] // U+5ABF <cjk>
	`嫚`: [u8(0xF2), 0x8A] // U+5ADA <cjk>
	`嫜`: [u8(0xF2), 0x8B] // U+5ADC <cjk>
	`嫠`: [u8(0xF2), 0x8C] // U+5AE0 <cjk>
	`嫥`: [u8(0xF2), 0x8D] // U+5AE5 <cjk>
	`嫰`: [u8(0xF2), 0x8E] // U+5AF0 <cjk>
	`嫮`: [u8(0xF2), 0x8F] // U+5AEE <cjk>
	`嫵`: [u8(0xF2), 0x90] // U+5AF5 <cjk>
	`嬀`: [u8(0xF2), 0x91] // U+5B00 <cjk>
	`嬈`: [u8(0xF2), 0x92] // U+5B08 <cjk>
	`嬗`: [u8(0xF2), 0x93] // U+5B17 <cjk>
	`嬴`: [u8(0xF2), 0x94] // U+5B34 <cjk>
	`嬭`: [u8(0xF2), 0x95] // U+5B2D <cjk>
	`孌`: [u8(0xF2), 0x96] // U+5B4C <cjk>
	`孒`: [u8(0xF2), 0x97] // U+5B52 <cjk>
	`孨`: [u8(0xF2), 0x98] // U+5B68 <cjk>
	`孯`: [u8(0xF2), 0x99] // U+5B6F <cjk>
	`孼`: [u8(0xF2), 0x9A] // U+5B7C <cjk>
	`孿`: [u8(0xF2), 0x9B] // U+5B7F <cjk>
	`宁`: [u8(0xF2), 0x9C] // U+5B81 <cjk>
	`宄`: [u8(0xF2), 0x9D] // U+5B84 <cjk>
	`𡧃`: [u8(0xF2), 0x9E] // U+219C3 <cjk>
	`幮`: [u8(0xF2), 0x9F] // U+5E6E <cjk>
	`𢅻`: [u8(0xF2), 0xA0] // U+2217B <cjk>
	`庥`: [u8(0xF2), 0xA1] // U+5EA5 <cjk>
	`庪`: [u8(0xF2), 0xA2] // U+5EAA <cjk>
	`庬`: [u8(0xF2), 0xA3] // U+5EAC <cjk>
	`庹`: [u8(0xF2), 0xA4] // U+5EB9 <cjk>
	`庿`: [u8(0xF2), 0xA5] // U+5EBF <cjk>
	`廆`: [u8(0xF2), 0xA6] // U+5EC6 <cjk>
	`廒`: [u8(0xF2), 0xA7] // U+5ED2 <cjk>
	`廙`: [u8(0xF2), 0xA8] // U+5ED9 <cjk>
	`𢌞`: [u8(0xF2), 0xA9] // U+2231E <cjk>
	`廽`: [u8(0xF2), 0xAA] // U+5EFD <cjk>
	`弈`: [u8(0xF2), 0xAB] // U+5F08 <cjk>
	`弎`: [u8(0xF2), 0xAC] // U+5F0E <cjk>
	`弜`: [u8(0xF2), 0xAD] // U+5F1C <cjk>
	`𢎭`: [u8(0xF2), 0xAE] // U+223AD <cjk>
	`弞`: [u8(0xF2), 0xAF] // U+5F1E <cjk>
	`彇`: [u8(0xF2), 0xB0] // U+5F47 <cjk>
	`彣`: [u8(0xF2), 0xB1] // U+5F63 <cjk>
	`彲`: [u8(0xF2), 0xB2] // U+5F72 <cjk>
	`彾`: [u8(0xF2), 0xB3] // U+5F7E <cjk>
	`徏`: [u8(0xF2), 0xB4] // U+5F8F <cjk>
	`徢`: [u8(0xF2), 0xB5] // U+5FA2 <cjk>
	`徤`: [u8(0xF2), 0xB6] // U+5FA4 <cjk>
	`徸`: [u8(0xF2), 0xB7] // U+5FB8 <cjk>
	`忄`: [u8(0xF2), 0xB8] // U+5FC4 <cjk>
	`㣺`: [u8(0xF2), 0xB9] // U+38FA <cjk>
	`忇`: [u8(0xF2), 0xBA] // U+5FC7 <cjk>
	`忋`: [u8(0xF2), 0xBB] // U+5FCB <cjk>
	`忒`: [u8(0xF2), 0xBC] // U+5FD2 <cjk>
	`忓`: [u8(0xF2), 0xBD] // U+5FD3 <cjk>
	`忔`: [u8(0xF2), 0xBE] // U+5FD4 <cjk>
	`忢`: [u8(0xF2), 0xBF] // U+5FE2 <cjk>
	`忮`: [u8(0xF2), 0xC0] // U+5FEE <cjk>
	`忯`: [u8(0xF2), 0xC1] // U+5FEF <cjk>
	`忳`: [u8(0xF2), 0xC2] // U+5FF3 <cjk>
	`忼`: [u8(0xF2), 0xC3] // U+5FFC <cjk>
	`㤗`: [u8(0xF2), 0xC4] // U+3917 <cjk>
	`怗`: [u8(0xF2), 0xC5] // U+6017 <cjk>
	`怢`: [u8(0xF2), 0xC6] // U+6022 <cjk>
	`怤`: [u8(0xF2), 0xC7] // U+6024 <cjk>
	`㤚`: [u8(0xF2), 0xC8] // U+391A <cjk>
	`恌`: [u8(0xF2), 0xC9] // U+604C <cjk>
	`恿`: [u8(0xF2), 0xCA] // U+607F <cjk>
	`悊`: [u8(0xF2), 0xCB] // U+608A <cjk>
	`悕`: [u8(0xF2), 0xCC] // U+6095 <cjk>
	`您`: [u8(0xF2), 0xCD] // U+60A8 <cjk>
	`𢛳`: [u8(0xF2), 0xCE] // U+226F3 <cjk>
	`悰`: [u8(0xF2), 0xCF] // U+60B0 <cjk>
	`悱`: [u8(0xF2), 0xD0] // U+60B1 <cjk>
	`悾`: [u8(0xF2), 0xD1] // U+60BE <cjk>
	`惈`: [u8(0xF2), 0xD2] // U+60C8 <cjk>
	`惙`: [u8(0xF2), 0xD3] // U+60D9 <cjk>
	`惛`: [u8(0xF2), 0xD4] // U+60DB <cjk>
	`惮`: [u8(0xF2), 0xD5] // U+60EE <cjk>
	`惲`: [u8(0xF2), 0xD6] // U+60F2 <cjk>
	`惵`: [u8(0xF2), 0xD7] // U+60F5 <cjk>
	`愐`: [u8(0xF2), 0xD8] // U+6110 <cjk>
	`愒`: [u8(0xF2), 0xD9] // U+6112 <cjk>
	`愓`: [u8(0xF2), 0xDA] // U+6113 <cjk>
	`愙`: [u8(0xF2), 0xDB] // U+6119 <cjk>
	`愞`: [u8(0xF2), 0xDC] // U+611E <cjk>
	`愺`: [u8(0xF2), 0xDD] // U+613A <cjk>
	`㥯`: [u8(0xF2), 0xDE] // U+396F <cjk>
	`慁`: [u8(0xF2), 0xDF] // U+6141 <cjk>
	`慆`: [u8(0xF2), 0xE0] // U+6146 <cjk>
	`慠`: [u8(0xF2), 0xE1] // U+6160 <cjk>
	`慼`: [u8(0xF2), 0xE2] // U+617C <cjk>
	`𢡛`: [u8(0xF2), 0xE3] // U+2285B <cjk>
	`憒`: [u8(0xF2), 0xE4] // U+6192 <cjk>
	`憓`: [u8(0xF2), 0xE5] // U+6193 <cjk>
	`憗`: [u8(0xF2), 0xE6] // U+6197 <cjk>
	`憘`: [u8(0xF2), 0xE7] // U+6198 <cjk>
	`憥`: [u8(0xF2), 0xE8] // U+61A5 <cjk>
	`憨`: [u8(0xF2), 0xE9] // U+61A8 <cjk>
	`憭`: [u8(0xF2), 0xEA] // U+61AD <cjk>
	`𢢫`: [u8(0xF2), 0xEB] // U+228AB <cjk>
	`懕`: [u8(0xF2), 0xEC] // U+61D5 <cjk>
	`懝`: [u8(0xF2), 0xED] // U+61DD <cjk>
	`懟`: [u8(0xF2), 0xEE] // U+61DF <cjk>
	`懵`: [u8(0xF2), 0xEF] // U+61F5 <cjk>
	`𢦏`: [u8(0xF2), 0xF0] // U+2298F <cjk>
	`戕`: [u8(0xF2), 0xF1] // U+6215 <cjk>
	`戣`: [u8(0xF2), 0xF2] // U+6223 <cjk>
	`戩`: [u8(0xF2), 0xF3] // U+6229 <cjk>
	`扆`: [u8(0xF2), 0xF4] // U+6246 <cjk>
	`扌`: [u8(0xF2), 0xF5] // U+624C <cjk>
	`扑`: [u8(0xF2), 0xF6] // U+6251 <cjk>
	`扒`: [u8(0xF2), 0xF7] // U+6252 <cjk>
	`扡`: [u8(0xF2), 0xF8] // U+6261 <cjk>
	`扤`: [u8(0xF2), 0xF9] // U+6264 <cjk>
	`扻`: [u8(0xF2), 0xFA] // U+627B <cjk>
	`扭`: [u8(0xF2), 0xFB] // U+626D <cjk>
	`扳`: [u8(0xF2), 0xFC] // U+6273 <cjk>
	`抙`: [u8(0xF3), 0x40] // U+6299 <cjk>
	`抦`: [u8(0xF3), 0x41] // U+62A6 <cjk>
	`拕`: [u8(0xF3), 0x42] // U+62D5 <cjk>
	`𢪸`: [u8(0xF3), 0x43] // U+22AB8 <cjk>
	`拽`: [u8(0xF3), 0x44] // U+62FD <cjk>
	`挃`: [u8(0xF3), 0x45] // U+6303 <cjk>
	`挍`: [u8(0xF3), 0x46] // U+630D <cjk>
	`挐`: [u8(0xF3), 0x47] // U+6310 <cjk>
	`𢭏`: [u8(0xF3), 0x48] // U+22B4F <cjk>
	`𢭐`: [u8(0xF3), 0x49] // U+22B50 <cjk>
	`挲`: [u8(0xF3), 0x4A] // U+6332 <cjk>
	`挵`: [u8(0xF3), 0x4B] // U+6335 <cjk>
	`挻`: [u8(0xF3), 0x4C] // U+633B <cjk>
	`挼`: [u8(0xF3), 0x4D] // U+633C <cjk>
	`捁`: [u8(0xF3), 0x4E] // U+6341 <cjk>
	`捄`: [u8(0xF3), 0x4F] // U+6344 <cjk>
	`捎`: [u8(0xF3), 0x50] // U+634E <cjk>
	`𢭆`: [u8(0xF3), 0x51] // U+22B46 <cjk>
	`捙`: [u8(0xF3), 0x52] // U+6359 <cjk>
	`𢰝`: [u8(0xF3), 0x53] // U+22C1D <cjk>
	`𢮦`: [u8(0xF3), 0x54] // U+22BA6 <cjk>
	`捬`: [u8(0xF3), 0x55] // U+636C <cjk>
	`掄`: [u8(0xF3), 0x56] // U+6384 <cjk>
	`掙`: [u8(0xF3), 0x57] // U+6399 <cjk>
	`𢰤`: [u8(0xF3), 0x58] // U+22C24 <cjk>
	`掔`: [u8(0xF3), 0x59] // U+6394 <cjk>
	`掽`: [u8(0xF3), 0x5A] // U+63BD <cjk>
	`揷`: [u8(0xF3), 0x5B] // U+63F7 <cjk>
	`揔`: [u8(0xF3), 0x5C] // U+63D4 <cjk>
	`揕`: [u8(0xF3), 0x5D] // U+63D5 <cjk>
	`揜`: [u8(0xF3), 0x5E] // U+63DC <cjk>
	`揠`: [u8(0xF3), 0x5F] // U+63E0 <cjk>
	`揫`: [u8(0xF3), 0x60] // U+63EB <cjk>
	`揬`: [u8(0xF3), 0x61] // U+63EC <cjk>
	`揲`: [u8(0xF3), 0x62] // U+63F2 <cjk>
	`搉`: [u8(0xF3), 0x63] // U+6409 <cjk>
	`搞`: [u8(0xF3), 0x64] // U+641E <cjk>
	`搥`: [u8(0xF3), 0x65] // U+6425 <cjk>
	`搩`: [u8(0xF3), 0x66] // U+6429 <cjk>
	`搯`: [u8(0xF3), 0x67] // U+642F <cjk>
	`摚`: [u8(0xF3), 0x68] // U+645A <cjk>
	`摛`: [u8(0xF3), 0x69] // U+645B <cjk>
	`摝`: [u8(0xF3), 0x6A] // U+645D <cjk>
	`摳`: [u8(0xF3), 0x6B] // U+6473 <cjk>
	`摽`: [u8(0xF3), 0x6C] // U+647D <cjk>
	`撇`: [u8(0xF3), 0x6D] // U+6487 <cjk>
	`撑`: [u8(0xF3), 0x6E] // U+6491 <cjk>
	`撝`: [u8(0xF3), 0x6F] // U+649D <cjk>
	`撟`: [u8(0xF3), 0x70] // U+649F <cjk>
	`擋`: [u8(0xF3), 0x71] // U+64CB <cjk>
	`擌`: [u8(0xF3), 0x72] // U+64CC <cjk>
	`擕`: [u8(0xF3), 0x73] // U+64D5 <cjk>
	`擗`: [u8(0xF3), 0x74] // U+64D7 <cjk>
	`𢷡`: [u8(0xF3), 0x75] // U+22DE1 <cjk>
	`擤`: [u8(0xF3), 0x76] // U+64E4 <cjk>
	`擥`: [u8(0xF3), 0x77] // U+64E5 <cjk>
	`擿`: [u8(0xF3), 0x78] // U+64FF <cjk>
	`攄`: [u8(0xF3), 0x79] // U+6504 <cjk>
	`㩮`: [u8(0xF3), 0x7A] // U+3A6E <cjk>
	`攏`: [u8(0xF3), 0x7B] // U+650F <cjk>
	`攔`: [u8(0xF3), 0x7C] // U+6514 <cjk>
	`攖`: [u8(0xF3), 0x7D] // U+6516 <cjk>
	`㩳`: [u8(0xF3), 0x7E] // U+3A73 <cjk>
	`攞`: [u8(0xF3), 0x80] // U+651E <cjk>
	`攲`: [u8(0xF3), 0x81] // U+6532 <cjk>
	`敄`: [u8(0xF3), 0x82] // U+6544 <cjk>
	`敔`: [u8(0xF3), 0x83] // U+6554 <cjk>
	`敫`: [u8(0xF3), 0x84] // U+656B <cjk>
	`敺`: [u8(0xF3), 0x85] // U+657A <cjk>
	`斁`: [u8(0xF3), 0x86] // U+6581 <cjk>
	`斄`: [u8(0xF3), 0x87] // U+6584 <cjk>
	`斅`: [u8(0xF3), 0x88] // U+6585 <cjk>
	`斊`: [u8(0xF3), 0x89] // U+658A <cjk>
	`斲`: [u8(0xF3), 0x8A] // U+65B2 <cjk>
	`斵`: [u8(0xF3), 0x8B] // U+65B5 <cjk>
	`斸`: [u8(0xF3), 0x8C] // U+65B8 <cjk>
	`斿`: [u8(0xF3), 0x8D] // U+65BF <cjk>
	`旂`: [u8(0xF3), 0x8E] // U+65C2 <cjk>
	`旉`: [u8(0xF3), 0x8F] // U+65C9 <cjk>
	`旔`: [u8(0xF3), 0x90] // U+65D4 <cjk>
	`㫖`: [u8(0xF3), 0x91] // U+3AD6 <cjk>
	`旲`: [u8(0xF3), 0x92] // U+65F2 <cjk>
	`旹`: [u8(0xF3), 0x93] // U+65F9 <cjk>
	`旼`: [u8(0xF3), 0x94] // U+65FC <cjk>
	`昄`: [u8(0xF3), 0x95] // U+6604 <cjk>
	`昈`: [u8(0xF3), 0x96] // U+6608 <cjk>
	`昡`: [u8(0xF3), 0x97] // U+6621 <cjk>
	`昪`: [u8(0xF3), 0x98] // U+662A <cjk>
	`晅`: [u8(0xF3), 0x99] // U+6645 <cjk>
	`晑`: [u8(0xF3), 0x9A] // U+6651 <cjk>
	`晎`: [u8(0xF3), 0x9B] // U+664E <cjk>
	`㫪`: [u8(0xF3), 0x9C] // U+3AEA <cjk>
	`𣇃`: [u8(0xF3), 0x9D] // U+231C3 <cjk>
	`晗`: [u8(0xF3), 0x9E] // U+6657 <cjk>
	`晛`: [u8(0xF3), 0x9F] // U+665B <cjk>
	`晣`: [u8(0xF3), 0xA0] // U+6663 <cjk>
	`𣇵`: [u8(0xF3), 0xA1] // U+231F5 <cjk>
	`𣆶`: [u8(0xF3), 0xA2] // U+231B6 <cjk>
	`晪`: [u8(0xF3), 0xA3] // U+666A <cjk>
	`晫`: [u8(0xF3), 0xA4] // U+666B <cjk>
	`晬`: [u8(0xF3), 0xA5] // U+666C <cjk>
	`晭`: [u8(0xF3), 0xA6] // U+666D <cjk>
	`晻`: [u8(0xF3), 0xA7] // U+667B <cjk>
	`暀`: [u8(0xF3), 0xA8] // U+6680 <cjk>
	`暐`: [u8(0xF3), 0xA9] // U+6690 <cjk>
	`暒`: [u8(0xF3), 0xAA] // U+6692 <cjk>
	`暙`: [u8(0xF3), 0xAB] // U+6699 <cjk>
	`㬎`: [u8(0xF3), 0xAC] // U+3B0E <cjk>
	`暭`: [u8(0xF3), 0xAD] // U+66AD <cjk>
	`暱`: [u8(0xF3), 0xAE] // U+66B1 <cjk>
	`暵`: [u8(0xF3), 0xAF] // U+66B5 <cjk>
	`㬚`: [u8(0xF3), 0xB0] // U+3B1A <cjk>
	`暿`: [u8(0xF3), 0xB1] // U+66BF <cjk>
	`㬜`: [u8(0xF3), 0xB2] // U+3B1C <cjk>
	`曬`: [u8(0xF3), 0xB3] // U+66EC <cjk>
	`㫗`: [u8(0xF3), 0xB4] // U+3AD7 <cjk>
	`朁`: [u8(0xF3), 0xB5] // U+6701 <cjk>
	`朅`: [u8(0xF3), 0xB6] // U+6705 <cjk>
	`朒`: [u8(0xF3), 0xB7] // U+6712 <cjk>
	`𣍲`: [u8(0xF3), 0xB8] // U+23372 <cjk>
	`朙`: [u8(0xF3), 0xB9] // U+6719 <cjk>
	`𣏓`: [u8(0xF3), 0xBA] // U+233D3 <cjk>
	`𣏒`: [u8(0xF3), 0xBB] // U+233D2 <cjk>
	`杌`: [u8(0xF3), 0xBC] // U+674C <cjk>
	`杍`: [u8(0xF3), 0xBD] // U+674D <cjk>
	`杔`: [u8(0xF3), 0xBE] // U+6754 <cjk>
	`杝`: [u8(0xF3), 0xBF] // U+675D <cjk>
	`𣏐`: [u8(0xF3), 0xC0] // U+233D0 <cjk>
	`𣏤`: [u8(0xF3), 0xC1] // U+233E4 <cjk>
	`𣏕`: [u8(0xF3), 0xC2] // U+233D5 <cjk>
	`杴`: [u8(0xF3), 0xC3] // U+6774 <cjk>
	`杶`: [u8(0xF3), 0xC4] // U+6776 <cjk>
	`𣏚`: [u8(0xF3), 0xC5] // U+233DA <cjk>
	`枒`: [u8(0xF3), 0xC6] // U+6792 <cjk>
	`𣏟`: [u8(0xF3), 0xC7] // U+233DF <cjk>
	`荣`: [u8(0xF3), 0xC8] // U+8363 <cjk>
	`栐`: [u8(0xF3), 0xC9] // U+6810 <cjk>
	`枰`: [u8(0xF3), 0xCA] // U+67B0 <cjk>
	`枲`: [u8(0xF3), 0xCB] // U+67B2 <cjk>
	`柃`: [u8(0xF3), 0xCC] // U+67C3 <cjk>
	`柈`: [u8(0xF3), 0xCD] // U+67C8 <cjk>
	`柒`: [u8(0xF3), 0xCE] // U+67D2 <cjk>
	`柙`: [u8(0xF3), 0xCF] // U+67D9 <cjk>
	`柛`: [u8(0xF3), 0xD0] // U+67DB <cjk>
	`柰`: [u8(0xF3), 0xD1] // U+67F0 <cjk>
	`柷`: [u8(0xF3), 0xD2] // U+67F7 <cjk>
	`𣑊`: [u8(0xF3), 0xD3] // U+2344A <cjk>
	`𣑑`: [u8(0xF3), 0xD4] // U+23451 <cjk>
	`𣑋`: [u8(0xF3), 0xD5] // U+2344B <cjk>
	`栘`: [u8(0xF3), 0xD6] // U+6818 <cjk>
	`栟`: [u8(0xF3), 0xD7] // U+681F <cjk>
	`栭`: [u8(0xF3), 0xD8] // U+682D <cjk>
	`𣑥`: [u8(0xF3), 0xD9] // U+23465 <cjk>
	`栳`: [u8(0xF3), 0xDA] // U+6833 <cjk>
	`栻`: [u8(0xF3), 0xDB] // U+683B <cjk>
	`栾`: [u8(0xF3), 0xDC] // U+683E <cjk>
	`桄`: [u8(0xF3), 0xDD] // U+6844 <cjk>
	`桅`: [u8(0xF3), 0xDE] // U+6845 <cjk>
	`桉`: [u8(0xF3), 0xDF] // U+6849 <cjk>
	`桌`: [u8(0xF3), 0xE0] // U+684C <cjk>
	`桕`: [u8(0xF3), 0xE1] // U+6855 <cjk>
	`桗`: [u8(0xF3), 0xE2] // U+6857 <cjk>
	`㭷`: [u8(0xF3), 0xE3] // U+3B77 <cjk>
	`桫`: [u8(0xF3), 0xE4] // U+686B <cjk>
	`桮`: [u8(0xF3), 0xE5] // U+686E <cjk>
	`桺`: [u8(0xF3), 0xE6] // U+687A <cjk>
	`桼`: [u8(0xF3), 0xE7] // U+687C <cjk>
	`梂`: [u8(0xF3), 0xE8] // U+6882 <cjk>
	`梐`: [u8(0xF3), 0xE9] // U+6890 <cjk>
	`梖`: [u8(0xF3), 0xEA] // U+6896 <cjk>
	`㭭`: [u8(0xF3), 0xEB] // U+3B6D <cjk>
	`梘`: [u8(0xF3), 0xEC] // U+6898 <cjk>
	`梙`: [u8(0xF3), 0xED] // U+6899 <cjk>
	`梚`: [u8(0xF3), 0xEE] // U+689A <cjk>
	`梜`: [u8(0xF3), 0xEF] // U+689C <cjk>
	`梪`: [u8(0xF3), 0xF0] // U+68AA <cjk>
	`梫`: [u8(0xF3), 0xF1] // U+68AB <cjk>
	`梴`: [u8(0xF3), 0xF2] // U+68B4 <cjk>
	`梻`: [u8(0xF3), 0xF3] // U+68BB <cjk>
	`棻`: [u8(0xF3), 0xF4] // U+68FB <cjk>
	`𣓤`: [u8(0xF3), 0xF5] // U+234E4 <cjk>
	`𣕚`: [u8(0xF3), 0xF6] // U+2355A <cjk>
	`﨓`: [u8(0xF3), 0xF7] // U+FA13 CJK COMPATIBILITY IDEOGRAPH-FA13
	`棃`: [u8(0xF3), 0xF8] // U+68C3 <cjk>
	`棅`: [u8(0xF3), 0xF9] // U+68C5 <cjk>
	`棌`: [u8(0xF3), 0xFA] // U+68CC <cjk>
	`棏`: [u8(0xF3), 0xFB] // U+68CF <cjk>
	`棖`: [u8(0xF3), 0xFC] // U+68D6 <cjk>
	`棙`: [u8(0xF4), 0x40] // U+68D9 <cjk>
	`棤`: [u8(0xF4), 0x41] // U+68E4 <cjk>
	`棥`: [u8(0xF4), 0x42] // U+68E5 <cjk>
	`棬`: [u8(0xF4), 0x43] // U+68EC <cjk>
	`棷`: [u8(0xF4), 0x44] // U+68F7 <cjk>
	`椃`: [u8(0xF4), 0x45] // U+6903 <cjk>
	`椇`: [u8(0xF4), 0x46] // U+6907 <cjk>
	`㮇`: [u8(0xF4), 0x47] // U+3B87 <cjk>
	`㮈`: [u8(0xF4), 0x48] // U+3B88 <cjk>
	`𣖔`: [u8(0xF4), 0x49] // U+23594 <cjk>
	`椻`: [u8(0xF4), 0x4A] // U+693B <cjk>
	`㮍`: [u8(0xF4), 0x4B] // U+3B8D <cjk>
	`楆`: [u8(0xF4), 0x4C] // U+6946 <cjk>
	`楩`: [u8(0xF4), 0x4D] // U+6969 <cjk>
	`楬`: [u8(0xF4), 0x4E] // U+696C <cjk>
	`楲`: [u8(0xF4), 0x4F] // U+6972 <cjk>
	`楺`: [u8(0xF4), 0x50] // U+697A <cjk>
	`楿`: [u8(0xF4), 0x51] // U+697F <cjk>
	`榒`: [u8(0xF4), 0x52] // U+6992 <cjk>
	`㮤`: [u8(0xF4), 0x53] // U+3BA4 <cjk>
	`榖`: [u8(0xF4), 0x54] // U+6996 <cjk>
	`榘`: [u8(0xF4), 0x55] // U+6998 <cjk>
	`榦`: [u8(0xF4), 0x56] // U+69A6 <cjk>
	`榰`: [u8(0xF4), 0x57] // U+69B0 <cjk>
	`榷`: [u8(0xF4), 0x58] // U+69B7 <cjk>
	`榺`: [u8(0xF4), 0x59] // U+69BA <cjk>
	`榼`: [u8(0xF4), 0x5A] // U+69BC <cjk>
	`槀`: [u8(0xF4), 0x5B] // U+69C0 <cjk>
	`槑`: [u8(0xF4), 0x5C] // U+69D1 <cjk>
	`槖`: [u8(0xF4), 0x5D] // U+69D6 <cjk>
	`𣘹`: [u8(0xF4), 0x5E] // U+23639 <cjk>
	`𣙇`: [u8(0xF4), 0x5F] // U+23647 <cjk>
	`樰`: [u8(0xF4), 0x60] // U+6A30 <cjk>
	`𣘸`: [u8(0xF4), 0x61] // U+23638 <cjk>
	`𣘺`: [u8(0xF4), 0x62] // U+2363A <cjk>
	`槣`: [u8(0xF4), 0x63] // U+69E3 <cjk>
	`槮`: [u8(0xF4), 0x64] // U+69EE <cjk>
	`槯`: [u8(0xF4), 0x65] // U+69EF <cjk>
	`槳`: [u8(0xF4), 0x66] // U+69F3 <cjk>
	`㯍`: [u8(0xF4), 0x67] // U+3BCD <cjk>
	`槴`: [u8(0xF4), 0x68] // U+69F4 <cjk>
	`槾`: [u8(0xF4), 0x69] // U+69FE <cjk>
	`樑`: [u8(0xF4), 0x6A] // U+6A11 <cjk>
	`樚`: [u8(0xF4), 0x6B] // U+6A1A <cjk>
	`樝`: [u8(0xF4), 0x6C] // U+6A1D <cjk>
	`𣜜`: [u8(0xF4), 0x6D] // U+2371C <cjk>
	`樲`: [u8(0xF4), 0x6E] // U+6A32 <cjk>
	`樳`: [u8(0xF4), 0x6F] // U+6A33 <cjk>
	`樴`: [u8(0xF4), 0x70] // U+6A34 <cjk>
	`樿`: [u8(0xF4), 0x71] // U+6A3F <cjk>
	`橆`: [u8(0xF4), 0x72] // U+6A46 <cjk>
	`橉`: [u8(0xF4), 0x73] // U+6A49 <cjk>
	`橺`: [u8(0xF4), 0x74] // U+6A7A <cjk>
	`橎`: [u8(0xF4), 0x75] // U+6A4E <cjk>
	`橒`: [u8(0xF4), 0x76] // U+6A52 <cjk>
	`橤`: [u8(0xF4), 0x77] // U+6A64 <cjk>
	`𣜌`: [u8(0xF4), 0x78] // U+2370C <cjk>
	`橾`: [u8(0xF4), 0x79] // U+6A7E <cjk>
	`檃`: [u8(0xF4), 0x7A] // U+6A83 <cjk>
	`檋`: [u8(0xF4), 0x7B] // U+6A8B <cjk>
	`㯰`: [u8(0xF4), 0x7C] // U+3BF0 <cjk>
	`檑`: [u8(0xF4), 0x7D] // U+6A91 <cjk>
	`檟`: [u8(0xF4), 0x7E] // U+6A9F <cjk>
	`檡`: [u8(0xF4), 0x80] // U+6AA1 <cjk>
	`𣝤`: [u8(0xF4), 0x81] // U+23764 <cjk>
	`檫`: [u8(0xF4), 0x82] // U+6AAB <cjk>
	`檽`: [u8(0xF4), 0x83] // U+6ABD <cjk>
	`櫆`: [u8(0xF4), 0x84] // U+6AC6 <cjk>
	`櫔`: [u8(0xF4), 0x85] // U+6AD4 <cjk>
	`櫐`: [u8(0xF4), 0x86] // U+6AD0 <cjk>
	`櫜`: [u8(0xF4), 0x87] // U+6ADC <cjk>
	`櫝`: [u8(0xF4), 0x88] // U+6ADD <cjk>
	`𣟿`: [u8(0xF4), 0x89] // U+237FF <cjk>
	`𣟧`: [u8(0xF4), 0x8A] // U+237E7 <cjk>
	`櫬`: [u8(0xF4), 0x8B] // U+6AEC <cjk>
	`櫱`: [u8(0xF4), 0x8C] // U+6AF1 <cjk>
	`櫲`: [u8(0xF4), 0x8D] // U+6AF2 <cjk>
	`櫳`: [u8(0xF4), 0x8E] // U+6AF3 <cjk>
	`櫽`: [u8(0xF4), 0x8F] // U+6AFD <cjk>
	`𣠤`: [u8(0xF4), 0x90] // U+23824 <cjk>
	`欋`: [u8(0xF4), 0x91] // U+6B0B <cjk>
	`欏`: [u8(0xF4), 0x92] // U+6B0F <cjk>
	`欐`: [u8(0xF4), 0x93] // U+6B10 <cjk>
	`欑`: [u8(0xF4), 0x94] // U+6B11 <cjk>
	`𣠽`: [u8(0xF4), 0x95] // U+2383D <cjk>
	`欗`: [u8(0xF4), 0x96] // U+6B17 <cjk>
	`㰦`: [u8(0xF4), 0x97] // U+3C26 <cjk>
	`欯`: [u8(0xF4), 0x98] // U+6B2F <cjk>
	`歊`: [u8(0xF4), 0x99] // U+6B4A <cjk>
	`歘`: [u8(0xF4), 0x9A] // U+6B58 <cjk>
	`歬`: [u8(0xF4), 0x9B] // U+6B6C <cjk>
	`歵`: [u8(0xF4), 0x9C] // U+6B75 <cjk>
	`歺`: [u8(0xF4), 0x9D] // U+6B7A <cjk>
	`殁`: [u8(0xF4), 0x9E] // U+6B81 <cjk>
	`殛`: [u8(0xF4), 0x9F] // U+6B9B <cjk>
	`殮`: [u8(0xF4), 0xA0] // U+6BAE <cjk>
	`𣪘`: [u8(0xF4), 0xA1] // U+23A98 <cjk>
	`殽`: [u8(0xF4), 0xA2] // U+6BBD <cjk>
	`殾`: [u8(0xF4), 0xA3] // U+6BBE <cjk>
	`毇`: [u8(0xF4), 0xA4] // U+6BC7 <cjk>
	`毈`: [u8(0xF4), 0xA5] // U+6BC8 <cjk>
	`毉`: [u8(0xF4), 0xA6] // U+6BC9 <cjk>
	`毚`: [u8(0xF4), 0xA7] // U+6BDA <cjk>
	`毦`: [u8(0xF4), 0xA8] // U+6BE6 <cjk>
	`毧`: [u8(0xF4), 0xA9] // U+6BE7 <cjk>
	`毮`: [u8(0xF4), 0xAA] // U+6BEE <cjk>
	`毱`: [u8(0xF4), 0xAB] // U+6BF1 <cjk>
	`氂`: [u8(0xF4), 0xAC] // U+6C02 <cjk>
	`氊`: [u8(0xF4), 0xAD] // U+6C0A <cjk>
	`氎`: [u8(0xF4), 0xAE] // U+6C0E <cjk>
	`氵`: [u8(0xF4), 0xAF] // U+6C35 <cjk>
	`氶`: [u8(0xF4), 0xB0] // U+6C36 <cjk>
	`氺`: [u8(0xF4), 0xB1] // U+6C3A <cjk>
	`𣱿`: [u8(0xF4), 0xB2] // U+23C7F <cjk>
	`氿`: [u8(0xF4), 0xB3] // U+6C3F <cjk>
	`汍`: [u8(0xF4), 0xB4] // U+6C4D <cjk>
	`汛`: [u8(0xF4), 0xB5] // U+6C5B <cjk>
	`汭`: [u8(0xF4), 0xB6] // U+6C6D <cjk>
	`沄`: [u8(0xF4), 0xB7] // U+6C84 <cjk>
	`沉`: [u8(0xF4), 0xB8] // U+6C89 <cjk>
	`㳃`: [u8(0xF4), 0xB9] // U+3CC3 <cjk>
	`沔`: [u8(0xF4), 0xBA] // U+6C94 <cjk>
	`沕`: [u8(0xF4), 0xBB] // U+6C95 <cjk>
	`沗`: [u8(0xF4), 0xBC] // U+6C97 <cjk>
	`沭`: [u8(0xF4), 0xBD] // U+6CAD <cjk>
	`泂`: [u8(0xF4), 0xBE] // U+6CC2 <cjk>
	`泐`: [u8(0xF4), 0xBF] // U+6CD0 <cjk>
	`㳒`: [u8(0xF4), 0xC0] // U+3CD2 <cjk>
	`泖`: [u8(0xF4), 0xC1] // U+6CD6 <cjk>
	`泚`: [u8(0xF4), 0xC2] // U+6CDA <cjk>
	`泜`: [u8(0xF4), 0xC3] // U+6CDC <cjk>
	`泩`: [u8(0xF4), 0xC4] // U+6CE9 <cjk>
	`泬`: [u8(0xF4), 0xC5] // U+6CEC <cjk>
	`泭`: [u8(0xF4), 0xC6] // U+6CED <cjk>
	`𣴀`: [u8(0xF4), 0xC7] // U+23D00 <cjk>
	`洀`: [u8(0xF4), 0xC8] // U+6D00 <cjk>
	`洊`: [u8(0xF4), 0xC9] // U+6D0A <cjk>
	`洤`: [u8(0xF4), 0xCA] // U+6D24 <cjk>
	`洦`: [u8(0xF4), 0xCB] // U+6D26 <cjk>
	`洧`: [u8(0xF4), 0xCC] // U+6D27 <cjk>
	`汧`: [u8(0xF4), 0xCD] // U+6C67 <cjk>
	`洯`: [u8(0xF4), 0xCE] // U+6D2F <cjk>
	`洼`: [u8(0xF4), 0xCF] // U+6D3C <cjk>
	`浛`: [u8(0xF4), 0xD0] // U+6D5B <cjk>
	`浞`: [u8(0xF4), 0xD1] // U+6D5E <cjk>
	`浠`: [u8(0xF4), 0xD2] // U+6D60 <cjk>
	`浰`: [u8(0xF4), 0xD3] // U+6D70 <cjk>
	`涀`: [u8(0xF4), 0xD4] // U+6D80 <cjk>
	`涁`: [u8(0xF4), 0xD5] // U+6D81 <cjk>
	`涊`: [u8(0xF4), 0xD6] // U+6D8A <cjk>
	`涍`: [u8(0xF4), 0xD7] // U+6D8D <cjk>
	`涑`: [u8(0xF4), 0xD8] // U+6D91 <cjk>
	`涘`: [u8(0xF4), 0xD9] // U+6D98 <cjk>
	`𣵀`: [u8(0xF4), 0xDA] // U+23D40 <cjk>
	`渗`: [u8(0xF4), 0xDB] // U+6E17 <cjk>
	`𣷺`: [u8(0xF4), 0xDC] // U+23DFA <cjk>
	`𣷹`: [u8(0xF4), 0xDD] // U+23DF9 <cjk>
	`𣷓`: [u8(0xF4), 0xDE] // U+23DD3 <cjk>
	`涫`: [u8(0xF4), 0xDF] // U+6DAB <cjk>
	`涮`: [u8(0xF4), 0xE0] // U+6DAE <cjk>
	`涴`: [u8(0xF4), 0xE1] // U+6DB4 <cjk>
	`淂`: [u8(0xF4), 0xE2] // U+6DC2 <cjk>
	`洴`: [u8(0xF4), 0xE3] // U+6D34 <cjk>
	`淈`: [u8(0xF4), 0xE4] // U+6DC8 <cjk>
	`淎`: [u8(0xF4), 0xE5] // U+6DCE <cjk>
	`淏`: [u8(0xF4), 0xE6] // U+6DCF <cjk>
	`淐`: [u8(0xF4), 0xE7] // U+6DD0 <cjk>
	`淟`: [u8(0xF4), 0xE8] // U+6DDF <cjk>
	`淩`: [u8(0xF4), 0xE9] // U+6DE9 <cjk>
	`淶`: [u8(0xF4), 0xEA] // U+6DF6 <cjk>
	`渶`: [u8(0xF4), 0xEB] // U+6E36 <cjk>
	`渞`: [u8(0xF4), 0xEC] // U+6E1E <cjk>
	`渢`: [u8(0xF4), 0xED] // U+6E22 <cjk>
	`渧`: [u8(0xF4), 0xEE] // U+6E27 <cjk>
	`㴑`: [u8(0xF4), 0xEF] // U+3D11 <cjk>
	`渲`: [u8(0xF4), 0xF0] // U+6E32 <cjk>
	`渼`: [u8(0xF4), 0xF1] // U+6E3C <cjk>
	`湈`: [u8(0xF4), 0xF2] // U+6E48 <cjk>
	`湉`: [u8(0xF4), 0xF3] // U+6E49 <cjk>
	`湋`: [u8(0xF4), 0xF4] // U+6E4B <cjk>
	`湌`: [u8(0xF4), 0xF5] // U+6E4C <cjk>
	`湏`: [u8(0xF4), 0xF6] // U+6E4F <cjk>
	`湑`: [u8(0xF4), 0xF7] // U+6E51 <cjk>
	`湓`: [u8(0xF4), 0xF8] // U+6E53 <cjk>
	`湔`: [u8(0xF4), 0xF9] // U+6E54 <cjk>
	`湗`: [u8(0xF4), 0xFA] // U+6E57 <cjk>
	`湣`: [u8(0xF4), 0xFB] // U+6E63 <cjk>
	`㴞`: [u8(0xF4), 0xFC] // U+3D1E <cjk>
	`溓`: [u8(0xF5), 0x40] // U+6E93 <cjk>
	`溧`: [u8(0xF5), 0x41] // U+6EA7 <cjk>
	`溴`: [u8(0xF5), 0x42] // U+6EB4 <cjk>
	`溿`: [u8(0xF5), 0x43] // U+6EBF <cjk>
	`滃`: [u8(0xF5), 0x44] // U+6EC3 <cjk>
	`滊`: [u8(0xF5), 0x45] // U+6ECA <cjk>
	`滙`: [u8(0xF5), 0x46] // U+6ED9 <cjk>
	`漵`: [u8(0xF5), 0x47] // U+6F35 <cjk>
	`滫`: [u8(0xF5), 0x48] // U+6EEB <cjk>
	`滹`: [u8(0xF5), 0x49] // U+6EF9 <cjk>
	`滻`: [u8(0xF5), 0x4A] // U+6EFB <cjk>
	`漊`: [u8(0xF5), 0x4B] // U+6F0A <cjk>
	`漌`: [u8(0xF5), 0x4C] // U+6F0C <cjk>
	`漘`: [u8(0xF5), 0x4D] // U+6F18 <cjk>
	`漥`: [u8(0xF5), 0x4E] // U+6F25 <cjk>
	`漶`: [u8(0xF5), 0x4F] // U+6F36 <cjk>
	`漼`: [u8(0xF5), 0x50] // U+6F3C <cjk>
	`𣽾`: [u8(0xF5), 0x51] // U+23F7E <cjk>
	`潒`: [u8(0xF5), 0x52] // U+6F52 <cjk>
	`潗`: [u8(0xF5), 0x53] // U+6F57 <cjk>
	`潚`: [u8(0xF5), 0x54] // U+6F5A <cjk>
	`潠`: [u8(0xF5), 0x55] // U+6F60 <cjk>
	`潨`: [u8(0xF5), 0x56] // U+6F68 <cjk>
	`澘`: [u8(0xF5), 0x57] // U+6F98 <cjk>
	`潽`: [u8(0xF5), 0x58] // U+6F7D <cjk>
	`澐`: [u8(0xF5), 0x59] // U+6F90 <cjk>
	`澖`: [u8(0xF5), 0x5A] // U+6F96 <cjk>
	`澾`: [u8(0xF5), 0x5B] // U+6FBE <cjk>
	`澟`: [u8(0xF5), 0x5C] // U+6F9F <cjk>
	`澥`: [u8(0xF5), 0x5D] // U+6FA5 <cjk>
	`澯`: [u8(0xF5), 0x5E] // U+6FAF <cjk>
	`㵤`: [u8(0xF5), 0x5F] // U+3D64 <cjk>
	`澵`: [u8(0xF5), 0x60] // U+6FB5 <cjk>
	`濈`: [u8(0xF5), 0x61] // U+6FC8 <cjk>
	`濉`: [u8(0xF5), 0x62] // U+6FC9 <cjk>
	`濚`: [u8(0xF5), 0x63] // U+6FDA <cjk>
	`濞`: [u8(0xF5), 0x64] // U+6FDE <cjk>
	`濩`: [u8(0xF5), 0x65] // U+6FE9 <cjk>
	`𤂖`: [u8(0xF5), 0x66] // U+24096 <cjk>
	`濼`: [u8(0xF5), 0x67] // U+6FFC <cjk>
	`瀀`: [u8(0xF5), 0x68] // U+7000 <cjk>
	`瀇`: [u8(0xF5), 0x69] // U+7007 <cjk>
	`瀊`: [u8(0xF5), 0x6A] // U+700A <cjk>
	`瀣`: [u8(0xF5), 0x6B] // U+7023 <cjk>
	`𤄃`: [u8(0xF5), 0x6C] // U+24103 <cjk>
	`瀹`: [u8(0xF5), 0x6D] // U+7039 <cjk>
	`瀺`: [u8(0xF5), 0x6E] // U+703A <cjk>
	`瀼`: [u8(0xF5), 0x6F] // U+703C <cjk>
	`灃`: [u8(0xF5), 0x70] // U+7043 <cjk>
	`灇`: [u8(0xF5), 0x71] // U+7047 <cjk>
	`灋`: [u8(0xF5), 0x72] // U+704B <cjk>
	`㶚`: [u8(0xF5), 0x73] // U+3D9A <cjk>
	`灔`: [u8(0xF5), 0x74] // U+7054 <cjk>
	`灥`: [u8(0xF5), 0x75] // U+7065 <cjk>
	`灩`: [u8(0xF5), 0x76] // U+7069 <cjk>
	`灬`: [u8(0xF5), 0x77] // U+706C <cjk>
	`灮`: [u8(0xF5), 0x78] // U+706E <cjk>
	`灶`: [u8(0xF5), 0x79] // U+7076 <cjk>
	`灾`: [u8(0xF5), 0x7A] // U+707E <cjk>
	`炁`: [u8(0xF5), 0x7B] // U+7081 <cjk>
	`炆`: [u8(0xF5), 0x7C] // U+7086 <cjk>
	`炕`: [u8(0xF5), 0x7D] // U+7095 <cjk>
	`炗`: [u8(0xF5), 0x7E] // U+7097 <cjk>
	`炻`: [u8(0xF5), 0x80] // U+70BB <cjk>
	`𤇆`: [u8(0xF5), 0x81] // U+241C6 <cjk>
	`炟`: [u8(0xF5), 0x82] // U+709F <cjk>
	`炱`: [u8(0xF5), 0x83] // U+70B1 <cjk>
	`𤇾`: [u8(0xF5), 0x84] // U+241FE <cjk>
	`烬`: [u8(0xF5), 0x85] // U+70EC <cjk>
	`烊`: [u8(0xF5), 0x86] // U+70CA <cjk>
	`烑`: [u8(0xF5), 0x87] // U+70D1 <cjk>
	`烓`: [u8(0xF5), 0x88] // U+70D3 <cjk>
	`烜`: [u8(0xF5), 0x89] // U+70DC <cjk>
	`焃`: [u8(0xF5), 0x8A] // U+7103 <cjk>
	`焄`: [u8(0xF5), 0x8B] // U+7104 <cjk>
	`焆`: [u8(0xF5), 0x8C] // U+7106 <cjk>
	`焇`: [u8(0xF5), 0x8D] // U+7107 <cjk>
	`焈`: [u8(0xF5), 0x8E] // U+7108 <cjk>
	`焌`: [u8(0xF5), 0x8F] // U+710C <cjk>
	`㷀`: [u8(0xF5), 0x90] // U+3DC0 <cjk>
	`焯`: [u8(0xF5), 0x91] // U+712F <cjk>
	`焱`: [u8(0xF5), 0x92] // U+7131 <cjk>
	`煐`: [u8(0xF5), 0x93] // U+7150 <cjk>
	`煊`: [u8(0xF5), 0x94] // U+714A <cjk>
	`煓`: [u8(0xF5), 0x95] // U+7153 <cjk>
	`煞`: [u8(0xF5), 0x96] // U+715E <cjk>
	`㷔`: [u8(0xF5), 0x97] // U+3DD4 <cjk>
	`熖`: [u8(0xF5), 0x98] // U+7196 <cjk>
	`熀`: [u8(0xF5), 0x99] // U+7180 <cjk>
	`熛`: [u8(0xF5), 0x9A] // U+719B <cjk>
	`熠`: [u8(0xF5), 0x9B] // U+71A0 <cjk>
	`熢`: [u8(0xF5), 0x9C] // U+71A2 <cjk>
	`熮`: [u8(0xF5), 0x9D] // U+71AE <cjk>
	`熯`: [u8(0xF5), 0x9E] // U+71AF <cjk>
	`熳`: [u8(0xF5), 0x9F] // U+71B3 <cjk>
	`𤎼`: [u8(0xF5), 0xA0] // U+243BC <cjk>
	`燋`: [u8(0xF5), 0xA1] // U+71CB <cjk>
	`燓`: [u8(0xF5), 0xA2] // U+71D3 <cjk>
	`燙`: [u8(0xF5), 0xA3] // U+71D9 <cjk>
	`燜`: [u8(0xF5), 0xA4] // U+71DC <cjk>
	`爇`: [u8(0xF5), 0xA5] // U+7207 <cjk>
	`㸅`: [u8(0xF5), 0xA6] // U+3E05 <cjk>
	`爫`: [u8(0xF5), 0xA7] // U+FA49 CJK COMPATIBILITY IDEOGRAPH-FA49
	`爫`: [u8(0xF5), 0xA8] // U+722B <cjk>
	`爴`: [u8(0xF5), 0xA9] // U+7234 <cjk>
	`爸`: [u8(0xF5), 0xAA] // U+7238 <cjk>
	`爹`: [u8(0xF5), 0xAB] // U+7239 <cjk>
	`丬`: [u8(0xF5), 0xAC] // U+4E2C <cjk>
	`牂`: [u8(0xF5), 0xAD] // U+7242 <cjk>
	`牓`: [u8(0xF5), 0xAE] // U+7253 <cjk>
	`牗`: [u8(0xF5), 0xAF] // U+7257 <cjk>
	`牣`: [u8(0xF5), 0xB0] // U+7263 <cjk>
	`𤘩`: [u8(0xF5), 0xB1] // U+24629 <cjk>
	`牮`: [u8(0xF5), 0xB2] // U+726E <cjk>
	`牯`: [u8(0xF5), 0xB3] // U+726F <cjk>
	`牸`: [u8(0xF5), 0xB4] // U+7278 <cjk>
	`牿`: [u8(0xF5), 0xB5] // U+727F <cjk>
	`犎`: [u8(0xF5), 0xB6] // U+728E <cjk>
	`𤚥`: [u8(0xF5), 0xB7] // U+246A5 <cjk>
	`犭`: [u8(0xF5), 0xB8] // U+72AD <cjk>
	`犮`: [u8(0xF5), 0xB9] // U+72AE <cjk>
	`犰`: [u8(0xF5), 0xBA] // U+72B0 <cjk>
	`犱`: [u8(0xF5), 0xBB] // U+72B1 <cjk>
	`狁`: [u8(0xF5), 0xBC] // U+72C1 <cjk>
	`㹠`: [u8(0xF5), 0xBD] // U+3E60 <cjk>
	`狌`: [u8(0xF5), 0xBE] // U+72CC <cjk>
	`㹦`: [u8(0xF5), 0xBF] // U+3E66 <cjk>
	`㹨`: [u8(0xF5), 0xC0] // U+3E68 <cjk>
	`狳`: [u8(0xF5), 0xC1] // U+72F3 <cjk>
	`狺`: [u8(0xF5), 0xC2] // U+72FA <cjk>
	`猇`: [u8(0xF5), 0xC3] // U+7307 <cjk>
	`猒`: [u8(0xF5), 0xC4] // U+7312 <cjk>
	`猘`: [u8(0xF5), 0xC5] // U+7318 <cjk>
	`猙`: [u8(0xF5), 0xC6] // U+7319 <cjk>
	`㺃`: [u8(0xF5), 0xC7] // U+3E83 <cjk>
	`猹`: [u8(0xF5), 0xC8] // U+7339 <cjk>
	`猬`: [u8(0xF5), 0xC9] // U+732C <cjk>
	`猱`: [u8(0xF5), 0xCA] // U+7331 <cjk>
	`猳`: [u8(0xF5), 0xCB] // U+7333 <cjk>
	`猽`: [u8(0xF5), 0xCC] // U+733D <cjk>
	`獒`: [u8(0xF5), 0xCD] // U+7352 <cjk>
	`㺔`: [u8(0xF5), 0xCE] // U+3E94 <cjk>
	`獫`: [u8(0xF5), 0xCF] // U+736B <cjk>
	`獬`: [u8(0xF5), 0xD0] // U+736C <cjk>
	`𤢖`: [u8(0xF5), 0xD1] // U+24896 <cjk>
	`獮`: [u8(0xF5), 0xD2] // U+736E <cjk>
	`獯`: [u8(0xF5), 0xD3] // U+736F <cjk>
	`獱`: [u8(0xF5), 0xD4] // U+7371 <cjk>
	`獷`: [u8(0xF5), 0xD5] // U+7377 <cjk>
	`玁`: [u8(0xF5), 0xD6] // U+7381 <cjk>
	`玅`: [u8(0xF5), 0xD7] // U+7385 <cjk>
	`玊`: [u8(0xF5), 0xD8] // U+738A <cjk>
	`玔`: [u8(0xF5), 0xD9] // U+7394 <cjk>
	`玘`: [u8(0xF5), 0xDA] // U+7398 <cjk>
	`玜`: [u8(0xF5), 0xDB] // U+739C <cjk>
	`玞`: [u8(0xF5), 0xDC] // U+739E <cjk>
	`玥`: [u8(0xF5), 0xDD] // U+73A5 <cjk>
	`玨`: [u8(0xF5), 0xDE] // U+73A8 <cjk>
	`玵`: [u8(0xF5), 0xDF] // U+73B5 <cjk>
	`玷`: [u8(0xF5), 0xE0] // U+73B7 <cjk>
	`玹`: [u8(0xF5), 0xE1] // U+73B9 <cjk>
	`玼`: [u8(0xF5), 0xE2] // U+73BC <cjk>
	`玿`: [u8(0xF5), 0xE3] // U+73BF <cjk>
	`珅`: [u8(0xF5), 0xE4] // U+73C5 <cjk>
	`珋`: [u8(0xF5), 0xE5] // U+73CB <cjk>
	`珡`: [u8(0xF5), 0xE6] // U+73E1 <cjk>
	`珧`: [u8(0xF5), 0xE7] // U+73E7 <cjk>
	`珹`: [u8(0xF5), 0xE8] // U+73F9 <cjk>
	`琓`: [u8(0xF5), 0xE9] // U+7413 <cjk>
	`珺`: [u8(0xF5), 0xEA] // U+73FA <cjk>
	`琁`: [u8(0xF5), 0xEB] // U+7401 <cjk>
	`琤`: [u8(0xF5), 0xEC] // U+7424 <cjk>
	`琱`: [u8(0xF5), 0xED] // U+7431 <cjk>
	`琹`: [u8(0xF5), 0xEE] // U+7439 <cjk>
	`瑓`: [u8(0xF5), 0xEF] // U+7453 <cjk>
	`瑀`: [u8(0xF5), 0xF0] // U+7440 <cjk>
	`瑃`: [u8(0xF5), 0xF1] // U+7443 <cjk>
	`瑍`: [u8(0xF5), 0xF2] // U+744D <cjk>
	`瑒`: [u8(0xF5), 0xF3] // U+7452 <cjk>
	`瑝`: [u8(0xF5), 0xF4] // U+745D <cjk>
	`瑱`: [u8(0xF5), 0xF5] // U+7471 <cjk>
	`璁`: [u8(0xF5), 0xF6] // U+7481 <cjk>
	`璅`: [u8(0xF5), 0xF7] // U+7485 <cjk>
	`璈`: [u8(0xF5), 0xF8] // U+7488 <cjk>
	`𤩍`: [u8(0xF5), 0xF9] // U+24A4D <cjk>
	`璒`: [u8(0xF5), 0xFA] // U+7492 <cjk>
	`璗`: [u8(0xF5), 0xFB] // U+7497 <cjk>
	`璙`: [u8(0xF5), 0xFC] // U+7499 <cjk>
	`璠`: [u8(0xF6), 0x40] // U+74A0 <cjk>
	`璡`: [u8(0xF6), 0x41] // U+74A1 <cjk>
	`璥`: [u8(0xF6), 0x42] // U+74A5 <cjk>
	`璪`: [u8(0xF6), 0x43] // U+74AA <cjk>
	`璫`: [u8(0xF6), 0x44] // U+74AB <cjk>
	`璹`: [u8(0xF6), 0x45] // U+74B9 <cjk>
	`璻`: [u8(0xF6), 0x46] // U+74BB <cjk>
	`璺`: [u8(0xF6), 0x47] // U+74BA <cjk>
	`瓖`: [u8(0xF6), 0x48] // U+74D6 <cjk>
	`瓘`: [u8(0xF6), 0x49] // U+74D8 <cjk>
	`瓞`: [u8(0xF6), 0x4A] // U+74DE <cjk>
	`瓯`: [u8(0xF6), 0x4B] // U+74EF <cjk>
	`瓫`: [u8(0xF6), 0x4C] // U+74EB <cjk>
	`𤭖`: [u8(0xF6), 0x4D] // U+24B56 <cjk>
	`瓺`: [u8(0xF6), 0x4E] // U+74FA <cjk>
	`𤭯`: [u8(0xF6), 0x4F] // U+24B6F <cjk>
	`甠`: [u8(0xF6), 0x50] // U+7520 <cjk>
	`甤`: [u8(0xF6), 0x51] // U+7524 <cjk>
	`甪`: [u8(0xF6), 0x52] // U+752A <cjk>
	`㽗`: [u8(0xF6), 0x53] // U+3F57 <cjk>
	`𤰖`: [u8(0xF6), 0x54] // U+24C16 <cjk>
	`甽`: [u8(0xF6), 0x55] // U+753D <cjk>
	`甾`: [u8(0xF6), 0x56] // U+753E <cjk>
	`畀`: [u8(0xF6), 0x57] // U+7540 <cjk>
	`畈`: [u8(0xF6), 0x58] // U+7548 <cjk>
	`畎`: [u8(0xF6), 0x59] // U+754E <cjk>
	`畐`: [u8(0xF6), 0x5A] // U+7550 <cjk>
	`畒`: [u8(0xF6), 0x5B] // U+7552 <cjk>
	`畬`: [u8(0xF6), 0x5C] // U+756C <cjk>
	`畲`: [u8(0xF6), 0x5D] // U+7572 <cjk>
	`畱`: [u8(0xF6), 0x5E] // U+7571 <cjk>
	`畺`: [u8(0xF6), 0x5F] // U+757A <cjk>
	`畽`: [u8(0xF6), 0x60] // U+757D <cjk>
	`畾`: [u8(0xF6), 0x61] // U+757E <cjk>
	`疁`: [u8(0xF6), 0x62] // U+7581 <cjk>
	`𤴔`: [u8(0xF6), 0x63] // U+24D14 <cjk>
	`疌`: [u8(0xF6), 0x64] // U+758C <cjk>
	`㽵`: [u8(0xF6), 0x65] // U+3F75 <cjk>
	`疢`: [u8(0xF6), 0x66] // U+75A2 <cjk>
	`㽷`: [u8(0xF6), 0x67] // U+3F77 <cjk>
	`疰`: [u8(0xF6), 0x68] // U+75B0 <cjk>
	`疷`: [u8(0xF6), 0x69] // U+75B7 <cjk>
	`疿`: [u8(0xF6), 0x6A] // U+75BF <cjk>
	`痀`: [u8(0xF6), 0x6B] // U+75C0 <cjk>
	`痆`: [u8(0xF6), 0x6C] // U+75C6 <cjk>
	`痏`: [u8(0xF6), 0x6D] // U+75CF <cjk>
	`痓`: [u8(0xF6), 0x6E] // U+75D3 <cjk>
	`痝`: [u8(0xF6), 0x6F] // U+75DD <cjk>
	`痟`: [u8(0xF6), 0x70] // U+75DF <cjk>
	`痠`: [u8(0xF6), 0x71] // U+75E0 <cjk>
	`痧`: [u8(0xF6), 0x72] // U+75E7 <cjk>
	`痬`: [u8(0xF6), 0x73] // U+75EC <cjk>
	`痮`: [u8(0xF6), 0x74] // U+75EE <cjk>
	`痱`: [u8(0xF6), 0x75] // U+75F1 <cjk>
	`痹`: [u8(0xF6), 0x76] // U+75F9 <cjk>
	`瘃`: [u8(0xF6), 0x77] // U+7603 <cjk>
	`瘘`: [u8(0xF6), 0x78] // U+7618 <cjk>
	`瘇`: [u8(0xF6), 0x79] // U+7607 <cjk>
	`瘏`: [u8(0xF6), 0x7A] // U+760F <cjk>
	`㾮`: [u8(0xF6), 0x7B] // U+3FAE <cjk>
	`𤸎`: [u8(0xF6), 0x7C] // U+24E0E <cjk>
	`瘓`: [u8(0xF6), 0x7D] // U+7613 <cjk>
	`瘛`: [u8(0xF6), 0x7E] // U+761B <cjk>
	`瘜`: [u8(0xF6), 0x80] // U+761C <cjk>
	`𤸷`: [u8(0xF6), 0x81] // U+24E37 <cjk>
	`瘥`: [u8(0xF6), 0x82] // U+7625 <cjk>
	`瘨`: [u8(0xF6), 0x83] // U+7628 <cjk>
	`瘼`: [u8(0xF6), 0x84] // U+763C <cjk>
	`瘳`: [u8(0xF6), 0x85] // U+7633 <cjk>
	`𤹪`: [u8(0xF6), 0x86] // U+24E6A <cjk>
	`㿉`: [u8(0xF6), 0x87] // U+3FC9 <cjk>
	`癁`: [u8(0xF6), 0x88] // U+7641 <cjk>
	`𤺋`: [u8(0xF6), 0x89] // U+24E8B <cjk>
	`癉`: [u8(0xF6), 0x8A] // U+7649 <cjk>
	`癕`: [u8(0xF6), 0x8B] // U+7655 <cjk>
	`㿗`: [u8(0xF6), 0x8C] // U+3FD7 <cjk>
	`癮`: [u8(0xF6), 0x8D] // U+766E <cjk>
	`皕`: [u8(0xF6), 0x8E] // U+7695 <cjk>
	`皜`: [u8(0xF6), 0x8F] // U+769C <cjk>
	`皡`: [u8(0xF6), 0x90] // U+76A1 <cjk>
	`皠`: [u8(0xF6), 0x91] // U+76A0 <cjk>
	`皧`: [u8(0xF6), 0x92] // U+76A7 <cjk>
	`皨`: [u8(0xF6), 0x93] // U+76A8 <cjk>
	`皯`: [u8(0xF6), 0x94] // U+76AF <cjk>
	`𥁊`: [u8(0xF6), 0x95] // U+2504A <cjk>
	`盉`: [u8(0xF6), 0x96] // U+76C9 <cjk>
	`𥁕`: [u8(0xF6), 0x97] // U+25055 <cjk>
	`盨`: [u8(0xF6), 0x98] // U+76E8 <cjk>
	`盬`: [u8(0xF6), 0x99] // U+76EC <cjk>
	`𥄢`: [u8(0xF6), 0x9A] // U+25122 <cjk>
	`眗`: [u8(0xF6), 0x9B] // U+7717 <cjk>
	`眚`: [u8(0xF6), 0x9C] // U+771A <cjk>
	`眭`: [u8(0xF6), 0x9D] // U+772D <cjk>
	`眵`: [u8(0xF6), 0x9E] // U+7735 <cjk>
	`𥆩`: [u8(0xF6), 0x9F] // U+251A9 <cjk>
	`䀹`: [u8(0xF6), 0xA0] // U+4039 <cjk>
	`𥇥`: [u8(0xF6), 0xA1] // U+251E5 <cjk>
	`𥇍`: [u8(0xF6), 0xA2] // U+251CD <cjk>
	`睘`: [u8(0xF6), 0xA3] // U+7758 <cjk>
	`睠`: [u8(0xF6), 0xA4] // U+7760 <cjk>
	`睪`: [u8(0xF6), 0xA5] // U+776A <cjk>
	`𥈞`: [u8(0xF6), 0xA6] // U+2521E <cjk>
	`睲`: [u8(0xF6), 0xA7] // U+7772 <cjk>
	`睼`: [u8(0xF6), 0xA8] // U+777C <cjk>
	`睽`: [u8(0xF6), 0xA9] // U+777D <cjk>
	`𥉌`: [u8(0xF6), 0xAA] // U+2524C <cjk>
	`䁘`: [u8(0xF6), 0xAB] // U+4058 <cjk>
	`瞚`: [u8(0xF6), 0xAC] // U+779A <cjk>
	`瞟`: [u8(0xF6), 0xAD] // U+779F <cjk>
	`瞢`: [u8(0xF6), 0xAE] // U+77A2 <cjk>
	`瞤`: [u8(0xF6), 0xAF] // U+77A4 <cjk>
	`瞩`: [u8(0xF6), 0xB0] // U+77A9 <cjk>
	`矞`: [u8(0xF6), 0xB1] // U+77DE <cjk>
	`矟`: [u8(0xF6), 0xB2] // U+77DF <cjk>
	`矤`: [u8(0xF6), 0xB3] // U+77E4 <cjk>
	`矦`: [u8(0xF6), 0xB4] // U+77E6 <cjk>
	`矪`: [u8(0xF6), 0xB5] // U+77EA <cjk>
	`矬`: [u8(0xF6), 0xB6] // U+77EC <cjk>
	`䂓`: [u8(0xF6), 0xB7] // U+4093 <cjk>
	`矰`: [u8(0xF6), 0xB8] // U+77F0 <cjk>
	`矴`: [u8(0xF6), 0xB9] // U+77F4 <cjk>
	`矻`: [u8(0xF6), 0xBA] // U+77FB <cjk>
	`𥐮`: [u8(0xF6), 0xBB] // U+2542E <cjk>
	`砅`: [u8(0xF6), 0xBC] // U+7805 <cjk>
	`砆`: [u8(0xF6), 0xBD] // U+7806 <cjk>
	`砉`: [u8(0xF6), 0xBE] // U+7809 <cjk>
	`砍`: [u8(0xF6), 0xBF] // U+780D <cjk>
	`砙`: [u8(0xF6), 0xC0] // U+7819 <cjk>
	`砡`: [u8(0xF6), 0xC1] // U+7821 <cjk>
	`砬`: [u8(0xF6), 0xC2] // U+782C <cjk>
	`硇`: [u8(0xF6), 0xC3] // U+7847 <cjk>
	`硤`: [u8(0xF6), 0xC4] // U+7864 <cjk>
	`硪`: [u8(0xF6), 0xC5] // U+786A <cjk>
	`𥓙`: [u8(0xF6), 0xC6] // U+254D9 <cjk>
	`碊`: [u8(0xF6), 0xC7] // U+788A <cjk>
	`碔`: [u8(0xF6), 0xC8] // U+7894 <cjk>
	`碤`: [u8(0xF6), 0xC9] // U+78A4 <cjk>
	`碝`: [u8(0xF6), 0xCA] // U+789D <cjk>
	`碞`: [u8(0xF6), 0xCB] // U+789E <cjk>
	`碟`: [u8(0xF6), 0xCC] // U+789F <cjk>
	`碻`: [u8(0xF6), 0xCD] // U+78BB <cjk>
	`磈`: [u8(0xF6), 0xCE] // U+78C8 <cjk>
	`磌`: [u8(0xF6), 0xCF] // U+78CC <cjk>
	`磎`: [u8(0xF6), 0xD0] // U+78CE <cjk>
	`磕`: [u8(0xF6), 0xD1] // U+78D5 <cjk>
	`磠`: [u8(0xF6), 0xD2] // U+78E0 <cjk>
	`磡`: [u8(0xF6), 0xD3] // U+78E1 <cjk>
	`磦`: [u8(0xF6), 0xD4] // U+78E6 <cjk>
	`磹`: [u8(0xF6), 0xD5] // U+78F9 <cjk>
	`磺`: [u8(0xF6), 0xD6] // U+78FA <cjk>
	`磻`: [u8(0xF6), 0xD7] // U+78FB <cjk>
	`磾`: [u8(0xF6), 0xD8] // U+78FE <cjk>
	`𥖧`: [u8(0xF6), 0xD9] // U+255A7 <cjk>
	`礐`: [u8(0xF6), 0xDA] // U+7910 <cjk>
	`礛`: [u8(0xF6), 0xDB] // U+791B <cjk>
	`礰`: [u8(0xF6), 0xDC] // U+7930 <cjk>
	`礥`: [u8(0xF6), 0xDD] // U+7925 <cjk>
	`礻`: [u8(0xF6), 0xDE] // U+793B <cjk>
	`祊`: [u8(0xF6), 0xDF] // U+794A <cjk>
	`祘`: [u8(0xF6), 0xE0] // U+7958 <cjk>
	`祛`: [u8(0xF6), 0xE1] // U+795B <cjk>
	`䄅`: [u8(0xF6), 0xE2] // U+4105 <cjk>
	`祧`: [u8(0xF6), 0xE3] // U+7967 <cjk>
	`祲`: [u8(0xF6), 0xE4] // U+7972 <cjk>
	`禔`: [u8(0xF6), 0xE5] // U+7994 <cjk>
	`禕`: [u8(0xF6), 0xE6] // U+7995 <cjk>
	`禖`: [u8(0xF6), 0xE7] // U+7996 <cjk>
	`禛`: [u8(0xF6), 0xE8] // U+799B <cjk>
	`禡`: [u8(0xF6), 0xE9] // U+79A1 <cjk>
	`禩`: [u8(0xF6), 0xEA] // U+79A9 <cjk>
	`禴`: [u8(0xF6), 0xEB] // U+79B4 <cjk>
	`离`: [u8(0xF6), 0xEC] // U+79BB <cjk>
	`秂`: [u8(0xF6), 0xED] // U+79C2 <cjk>
	`秇`: [u8(0xF6), 0xEE] // U+79C7 <cjk>
	`秌`: [u8(0xF6), 0xEF] // U+79CC <cjk>
	`种`: [u8(0xF6), 0xF0] // U+79CD <cjk>
	`秖`: [u8(0xF6), 0xF1] // U+79D6 <cjk>
	`䅈`: [u8(0xF6), 0xF2] // U+4148 <cjk>
	`𥞩`: [u8(0xF6), 0xF3] // U+257A9 <cjk>
	`𥞴`: [u8(0xF6), 0xF4] // U+257B4 <cjk>
	`䅏`: [u8(0xF6), 0xF5] // U+414F <cjk>
	`稊`: [u8(0xF6), 0xF6] // U+7A0A <cjk>
	`稑`: [u8(0xF6), 0xF7] // U+7A11 <cjk>
	`稕`: [u8(0xF6), 0xF8] // U+7A15 <cjk>
	`稛`: [u8(0xF6), 0xF9] // U+7A1B <cjk>
	`稞`: [u8(0xF6), 0xFA] // U+7A1E <cjk>
	`䅣`: [u8(0xF6), 0xFB] // U+4163 <cjk>
	`稭`: [u8(0xF6), 0xFC] // U+7A2D <cjk>
	`稸`: [u8(0xF7), 0x40] // U+7A38 <cjk>
	`穇`: [u8(0xF7), 0x41] // U+7A47 <cjk>
	`穌`: [u8(0xF7), 0x42] // U+7A4C <cjk>
	`穖`: [u8(0xF7), 0x43] // U+7A56 <cjk>
	`穙`: [u8(0xF7), 0x44] // U+7A59 <cjk>
	`穜`: [u8(0xF7), 0x45] // U+7A5C <cjk>
	`穟`: [u8(0xF7), 0x46] // U+7A5F <cjk>
	`穠`: [u8(0xF7), 0x47] // U+7A60 <cjk>
	`穧`: [u8(0xF7), 0x48] // U+7A67 <cjk>
	`穪`: [u8(0xF7), 0x49] // U+7A6A <cjk>
	`穵`: [u8(0xF7), 0x4A] // U+7A75 <cjk>
	`穸`: [u8(0xF7), 0x4B] // U+7A78 <cjk>
	`窂`: [u8(0xF7), 0x4C] // U+7A82 <cjk>
	`窊`: [u8(0xF7), 0x4D] // U+7A8A <cjk>
	`窐`: [u8(0xF7), 0x4E] // U+7A90 <cjk>
	`窣`: [u8(0xF7), 0x4F] // U+7AA3 <cjk>
	`窬`: [u8(0xF7), 0x50] // U+7AAC <cjk>
	`𥧔`: [u8(0xF7), 0x51] // U+259D4 <cjk>
	`䆴`: [u8(0xF7), 0x52] // U+41B4 <cjk>
	`窹`: [u8(0xF7), 0x53] // U+7AB9 <cjk>
	`窼`: [u8(0xF7), 0x54] // U+7ABC <cjk>
	`窾`: [u8(0xF7), 0x55] // U+7ABE <cjk>
	`䆿`: [u8(0xF7), 0x56] // U+41BF <cjk>
	`竌`: [u8(0xF7), 0x57] // U+7ACC <cjk>
	`竑`: [u8(0xF7), 0x58] // U+7AD1 <cjk>
	`竧`: [u8(0xF7), 0x59] // U+7AE7 <cjk>
	`竨`: [u8(0xF7), 0x5A] // U+7AE8 <cjk>
	`竴`: [u8(0xF7), 0x5B] // U+7AF4 <cjk>
	`𥫤`: [u8(0xF7), 0x5C] // U+25AE4 <cjk>
	`𥫣`: [u8(0xF7), 0x5D] // U+25AE3 <cjk>
	`笇`: [u8(0xF7), 0x5E] // U+7B07 <cjk>
	`𥫱`: [u8(0xF7), 0x5F] // U+25AF1 <cjk>
	`笽`: [u8(0xF7), 0x60] // U+7B3D <cjk>
	`笧`: [u8(0xF7), 0x61] // U+7B27 <cjk>
	`笪`: [u8(0xF7), 0x62] // U+7B2A <cjk>
	`笮`: [u8(0xF7), 0x63] // U+7B2E <cjk>
	`笯`: [u8(0xF7), 0x64] // U+7B2F <cjk>
	`笱`: [u8(0xF7), 0x65] // U+7B31 <cjk>
	`䇦`: [u8(0xF7), 0x66] // U+41E6 <cjk>
	`䇳`: [u8(0xF7), 0x67] // U+41F3 <cjk>
	`筿`: [u8(0xF7), 0x68] // U+7B7F <cjk>
	`筁`: [u8(0xF7), 0x69] // U+7B41 <cjk>
	`䇮`: [u8(0xF7), 0x6A] // U+41EE <cjk>
	`筕`: [u8(0xF7), 0x6B] // U+7B55 <cjk>
	`筹`: [u8(0xF7), 0x6C] // U+7B79 <cjk>
	`筤`: [u8(0xF7), 0x6D] // U+7B64 <cjk>
	`筦`: [u8(0xF7), 0x6E] // U+7B66 <cjk>
	`筩`: [u8(0xF7), 0x6F] // U+7B69 <cjk>
	`筳`: [u8(0xF7), 0x70] // U+7B73 <cjk>
	`𥮲`: [u8(0xF7), 0x71] // U+25BB2 <cjk>
	`䈇`: [u8(0xF7), 0x72] // U+4207 <cjk>
	`箐`: [u8(0xF7), 0x73] // U+7B90 <cjk>
	`箑`: [u8(0xF7), 0x74] // U+7B91 <cjk>
	`箛`: [u8(0xF7), 0x75] // U+7B9B <cjk>
	`䈎`: [u8(0xF7), 0x76] // U+420E <cjk>
	`箯`: [u8(0xF7), 0x77] // U+7BAF <cjk>
	`箵`: [u8(0xF7), 0x78] // U+7BB5 <cjk>
	`箼`: [u8(0xF7), 0x79] // U+7BBC <cjk>
	`篅`: [u8(0xF7), 0x7A] // U+7BC5 <cjk>
	`篊`: [u8(0xF7), 0x7B] // U+7BCA <cjk>
	`𥱋`: [u8(0xF7), 0x7C] // U+25C4B <cjk>
	`𥱤`: [u8(0xF7), 0x7D] // U+25C64 <cjk>
	`篔`: [u8(0xF7), 0x7E] // U+7BD4 <cjk>
	`篖`: [u8(0xF7), 0x80] // U+7BD6 <cjk>
	`篚`: [u8(0xF7), 0x81] // U+7BDA <cjk>
	`篪`: [u8(0xF7), 0x82] // U+7BEA <cjk>
	`篰`: [u8(0xF7), 0x83] // U+7BF0 <cjk>
	`簃`: [u8(0xF7), 0x84] // U+7C03 <cjk>
	`簋`: [u8(0xF7), 0x85] // U+7C0B <cjk>
	`簎`: [u8(0xF7), 0x86] // U+7C0E <cjk>
	`簏`: [u8(0xF7), 0x87] // U+7C0F <cjk>
	`簦`: [u8(0xF7), 0x88] // U+7C26 <cjk>
	`籅`: [u8(0xF7), 0x89] // U+7C45 <cjk>
	`籊`: [u8(0xF7), 0x8A] // U+7C4A <cjk>
	`籑`: [u8(0xF7), 0x8B] // U+7C51 <cjk>
	`籗`: [u8(0xF7), 0x8C] // U+7C57 <cjk>
	`籞`: [u8(0xF7), 0x8D] // U+7C5E <cjk>
	`籡`: [u8(0xF7), 0x8E] // U+7C61 <cjk>
	`籩`: [u8(0xF7), 0x8F] // U+7C69 <cjk>
	`籮`: [u8(0xF7), 0x90] // U+7C6E <cjk>
	`籯`: [u8(0xF7), 0x91] // U+7C6F <cjk>
	`籰`: [u8(0xF7), 0x92] // U+7C70 <cjk>
	`𥸮`: [u8(0xF7), 0x93] // U+25E2E <cjk>
	`𥹖`: [u8(0xF7), 0x94] // U+25E56 <cjk>
	`𥹥`: [u8(0xF7), 0x95] // U+25E65 <cjk>
	`粦`: [u8(0xF7), 0x96] // U+7CA6 <cjk>
	`𥹢`: [u8(0xF7), 0x97] // U+25E62 <cjk>
	`粶`: [u8(0xF7), 0x98] // U+7CB6 <cjk>
	`粷`: [u8(0xF7), 0x99] // U+7CB7 <cjk>
	`粿`: [u8(0xF7), 0x9A] // U+7CBF <cjk>
	`𥻘`: [u8(0xF7), 0x9B] // U+25ED8 <cjk>
	`糄`: [u8(0xF7), 0x9C] // U+7CC4 <cjk>
	`𥻂`: [u8(0xF7), 0x9D] // U+25EC2 <cjk>
	`糈`: [u8(0xF7), 0x9E] // U+7CC8 <cjk>
	`糍`: [u8(0xF7), 0x9F] // U+7CCD <cjk>
	`𥻨`: [u8(0xF7), 0xA0] // U+25EE8 <cjk>
	`糗`: [u8(0xF7), 0xA1] // U+7CD7 <cjk>
	`𥼣`: [u8(0xF7), 0xA2] // U+25F23 <cjk>
	`糦`: [u8(0xF7), 0xA3] // U+7CE6 <cjk>
	`糫`: [u8(0xF7), 0xA4] // U+7CEB <cjk>
	`𥽜`: [u8(0xF7), 0xA5] // U+25F5C <cjk>
	`糵`: [u8(0xF7), 0xA6] // U+7CF5 <cjk>
	`紃`: [u8(0xF7), 0xA7] // U+7D03 <cjk>
	`紉`: [u8(0xF7), 0xA8] // U+7D09 <cjk>
	`䋆`: [u8(0xF7), 0xA9] // U+42C6 <cjk>
	`紒`: [u8(0xF7), 0xAA] // U+7D12 <cjk>
	`紞`: [u8(0xF7), 0xAB] // U+7D1E <cjk>
	`𥿠`: [u8(0xF7), 0xAC] // U+25FE0 <cjk>
	`𥿔`: [u8(0xF7), 0xAD] // U+25FD4 <cjk>
	`紽`: [u8(0xF7), 0xAE] // U+7D3D <cjk>
	`紾`: [u8(0xF7), 0xAF] // U+7D3E <cjk>
	`絀`: [u8(0xF7), 0xB0] // U+7D40 <cjk>
	`絇`: [u8(0xF7), 0xB1] // U+7D47 <cjk>
	`𦀌`: [u8(0xF7), 0xB2] // U+2600C <cjk>
	`𥿻`: [u8(0xF7), 0xB3] // U+25FFB <cjk>
	`䋖`: [u8(0xF7), 0xB4] // U+42D6 <cjk>
	`絙`: [u8(0xF7), 0xB5] // U+7D59 <cjk>
	`絚`: [u8(0xF7), 0xB6] // U+7D5A <cjk>
	`絪`: [u8(0xF7), 0xB7] // U+7D6A <cjk>
	`絰`: [u8(0xF7), 0xB8] // U+7D70 <cjk>
	`䋝`: [u8(0xF7), 0xB9] // U+42DD <cjk>
	`絿`: [u8(0xF7), 0xBA] // U+7D7F <cjk>
	`𦀗`: [u8(0xF7), 0xBB] // U+26017 <cjk>
	`綆`: [u8(0xF7), 0xBC] // U+7D86 <cjk>
	`綈`: [u8(0xF7), 0xBD] // U+7D88 <cjk>
	`綌`: [u8(0xF7), 0xBE] // U+7D8C <cjk>
	`綗`: [u8(0xF7), 0xBF] // U+7D97 <cjk>
	`𦁠`: [u8(0xF7), 0xC0] // U+26060 <cjk>
	`綝`: [u8(0xF7), 0xC1] // U+7D9D <cjk>
	`綧`: [u8(0xF7), 0xC2] // U+7DA7 <cjk>
	`綪`: [u8(0xF7), 0xC3] // U+7DAA <cjk>
	`綶`: [u8(0xF7), 0xC4] // U+7DB6 <cjk>
	`綷`: [u8(0xF7), 0xC5] // U+7DB7 <cjk>
	`緀`: [u8(0xF7), 0xC6] // U+7DC0 <cjk>
	`緗`: [u8(0xF7), 0xC7] // U+7DD7 <cjk>
	`緙`: [u8(0xF7), 0xC8] // U+7DD9 <cjk>
	`緦`: [u8(0xF7), 0xC9] // U+7DE6 <cjk>
	`緱`: [u8(0xF7), 0xCA] // U+7DF1 <cjk>
	`緹`: [u8(0xF7), 0xCB] // U+7DF9 <cjk>
	`䌂`: [u8(0xF7), 0xCC] // U+4302 <cjk>
	`𦃭`: [u8(0xF7), 0xCD] // U+260ED <cjk>
	`縉`: [u8(0xF7), 0xCE] // U+FA58 CJK COMPATIBILITY IDEOGRAPH-FA58
	`縐`: [u8(0xF7), 0xCF] // U+7E10 <cjk>
	`縗`: [u8(0xF7), 0xD0] // U+7E17 <cjk>
	`縝`: [u8(0xF7), 0xD1] // U+7E1D <cjk>
	`縠`: [u8(0xF7), 0xD2] // U+7E20 <cjk>
	`縧`: [u8(0xF7), 0xD3] // U+7E27 <cjk>
	`縬`: [u8(0xF7), 0xD4] // U+7E2C <cjk>
	`繅`: [u8(0xF7), 0xD5] // U+7E45 <cjk>
	`繳`: [u8(0xF7), 0xD6] // U+7E73 <cjk>
	`繵`: [u8(0xF7), 0xD7] // U+7E75 <cjk>
	`繾`: [u8(0xF7), 0xD8] // U+7E7E <cjk>
	`纆`: [u8(0xF7), 0xD9] // U+7E86 <cjk>
	`纇`: [u8(0xF7), 0xDA] // U+7E87 <cjk>
	`䌫`: [u8(0xF7), 0xDB] // U+432B <cjk>
	`纑`: [u8(0xF7), 0xDC] // U+7E91 <cjk>
	`纘`: [u8(0xF7), 0xDD] // U+7E98 <cjk>
	`纚`: [u8(0xF7), 0xDE] // U+7E9A <cjk>
	`䍃`: [u8(0xF7), 0xDF] // U+4343 <cjk>
	`缼`: [u8(0xF7), 0xE0] // U+7F3C <cjk>
	`缻`: [u8(0xF7), 0xE1] // U+7F3B <cjk>
	`缾`: [u8(0xF7), 0xE2] // U+7F3E <cjk>
	`罃`: [u8(0xF7), 0xE3] // U+7F43 <cjk>
	`罄`: [u8(0xF7), 0xE4] // U+7F44 <cjk>
	`罏`: [u8(0xF7), 0xE5] // U+7F4F <cjk>
	`㓁`: [u8(0xF7), 0xE6] // U+34C1 <cjk>
	`𦉰`: [u8(0xF7), 0xE7] // U+26270 <cjk>
	`罒`: [u8(0xF7), 0xE8] // U+7F52 <cjk>
	`𦊆`: [u8(0xF7), 0xE9] // U+26286 <cjk>
	`罡`: [u8(0xF7), 0xEA] // U+7F61 <cjk>
	`罣`: [u8(0xF7), 0xEB] // U+7F63 <cjk>
	`罤`: [u8(0xF7), 0xEC] // U+7F64 <cjk>
	`罭`: [u8(0xF7), 0xED] // U+7F6D <cjk>
	`罽`: [u8(0xF7), 0xEE] // U+7F7D <cjk>
	`罾`: [u8(0xF7), 0xEF] // U+7F7E <cjk>
	`𦍌`: [u8(0xF7), 0xF0] // U+2634C <cjk>
	`羐`: [u8(0xF7), 0xF1] // U+7F90 <cjk>
	`养`: [u8(0xF7), 0xF2] // U+517B <cjk>
	`𣴎`: [u8(0xF7), 0xF3] // U+23D0E <cjk>
	`羖`: [u8(0xF7), 0xF4] // U+7F96 <cjk>
	`羜`: [u8(0xF7), 0xF5] // U+7F9C <cjk>
	`羭`: [u8(0xF7), 0xF6] // U+7FAD <cjk>
	`𦐂`: [u8(0xF7), 0xF7] // U+26402 <cjk>
	`翃`: [u8(0xF7), 0xF8] // U+7FC3 <cjk>
	`翏`: [u8(0xF7), 0xF9] // U+7FCF <cjk>
	`翣`: [u8(0xF7), 0xFA] // U+7FE3 <cjk>
	`翥`: [u8(0xF7), 0xFB] // U+7FE5 <cjk>
	`翯`: [u8(0xF7), 0xFC] // U+7FEF <cjk>
	`翲`: [u8(0xF8), 0x40] // U+7FF2 <cjk>
	`耂`: [u8(0xF8), 0x41] // U+8002 <cjk>
	`耊`: [u8(0xF8), 0x42] // U+800A <cjk>
	`耈`: [u8(0xF8), 0x43] // U+8008 <cjk>
	`耎`: [u8(0xF8), 0x44] // U+800E <cjk>
	`耑`: [u8(0xF8), 0x45] // U+8011 <cjk>
	`耖`: [u8(0xF8), 0x46] // U+8016 <cjk>
	`耤`: [u8(0xF8), 0x47] // U+8024 <cjk>
	`耬`: [u8(0xF8), 0x48] // U+802C <cjk>
	`耰`: [u8(0xF8), 0x49] // U+8030 <cjk>
	`聃`: [u8(0xF8), 0x4A] // U+8043 <cjk>
	`聦`: [u8(0xF8), 0x4B] // U+8066 <cjk>
	`聱`: [u8(0xF8), 0x4C] // U+8071 <cjk>
	`聵`: [u8(0xF8), 0x4D] // U+8075 <cjk>
	`聻`: [u8(0xF8), 0x4E] // U+807B <cjk>
	`肙`: [u8(0xF8), 0x4F] // U+8099 <cjk>
	`肜`: [u8(0xF8), 0x50] // U+809C <cjk>
	`肤`: [u8(0xF8), 0x51] // U+80A4 <cjk>
	`肧`: [u8(0xF8), 0x52] // U+80A7 <cjk>
	`肸`: [u8(0xF8), 0x53] // U+80B8 <cjk>
	`𦙾`: [u8(0xF8), 0x54] // U+2667E <cjk>
	`胅`: [u8(0xF8), 0x55] // U+80C5 <cjk>
	`胕`: [u8(0xF8), 0x56] // U+80D5 <cjk>
	`胘`: [u8(0xF8), 0x57] // U+80D8 <cjk>
	`胦`: [u8(0xF8), 0x58] // U+80E6 <cjk>
	`𦚰`: [u8(0xF8), 0x59] // U+266B0 <cjk>
	`脍`: [u8(0xF8), 0x5A] // U+810D <cjk>
	`胵`: [u8(0xF8), 0x5B] // U+80F5 <cjk>
	`胻`: [u8(0xF8), 0x5C] // U+80FB <cjk>
	`䏮`: [u8(0xF8), 0x5D] // U+43EE <cjk>
	`脵`: [u8(0xF8), 0x5E] // U+8135 <cjk>
	`脖`: [u8(0xF8), 0x5F] // U+8116 <cjk>
	`脞`: [u8(0xF8), 0x60] // U+811E <cjk>
	`䏰`: [u8(0xF8), 0x61] // U+43F0 <cjk>
	`脤`: [u8(0xF8), 0x62] // U+8124 <cjk>
	`脧`: [u8(0xF8), 0x63] // U+8127 <cjk>
	`脬`: [u8(0xF8), 0x64] // U+812C <cjk>
	`𦜝`: [u8(0xF8), 0x65] // U+2671D <cjk>
	`脽`: [u8(0xF8), 0x66] // U+813D <cjk>
	`䐈`: [u8(0xF8), 0x67] // U+4408 <cjk>
	`腩`: [u8(0xF8), 0x68] // U+8169 <cjk>
	`䐗`: [u8(0xF8), 0x69] // U+4417 <cjk>
	`膁`: [u8(0xF8), 0x6A] // U+8181 <cjk>
	`䐜`: [u8(0xF8), 0x6B] // U+441C <cjk>
	`膄`: [u8(0xF8), 0x6C] // U+8184 <cjk>
	`膅`: [u8(0xF8), 0x6D] // U+8185 <cjk>
	`䐢`: [u8(0xF8), 0x6E] // U+4422 <cjk>
	`膘`: [u8(0xF8), 0x6F] // U+8198 <cjk>
	`膲`: [u8(0xF8), 0x70] // U+81B2 <cjk>
	`臁`: [u8(0xF8), 0x71] // U+81C1 <cjk>
	`臃`: [u8(0xF8), 0x72] // U+81C3 <cjk>
	`臖`: [u8(0xF8), 0x73] // U+81D6 <cjk>
	`臛`: [u8(0xF8), 0x74] // U+81DB <cjk>
	`𦣝`: [u8(0xF8), 0x75] // U+268DD <cjk>
	`臤`: [u8(0xF8), 0x76] // U+81E4 <cjk>
	`𦣪`: [u8(0xF8), 0x77] // U+268EA <cjk>
	`臬`: [u8(0xF8), 0x78] // U+81EC <cjk>
	`𦥑`: [u8(0xF8), 0x79] // U+26951 <cjk>
	`臽`: [u8(0xF8), 0x7A] // U+81FD <cjk>
	`臿`: [u8(0xF8), 0x7B] // U+81FF <cjk>
	`𦥯`: [u8(0xF8), 0x7C] // U+2696F <cjk>
	`舄`: [u8(0xF8), 0x7D] // U+8204 <cjk>
	`𦧝`: [u8(0xF8), 0x7E] // U+269DD <cjk>
	`舙`: [u8(0xF8), 0x80] // U+8219 <cjk>
	`舡`: [u8(0xF8), 0x81] // U+8221 <cjk>
	`舢`: [u8(0xF8), 0x82] // U+8222 <cjk>
	`𦨞`: [u8(0xF8), 0x83] // U+26A1E <cjk>
	`舲`: [u8(0xF8), 0x84] // U+8232 <cjk>
	`舴`: [u8(0xF8), 0x85] // U+8234 <cjk>
	`舼`: [u8(0xF8), 0x86] // U+823C <cjk>
	`艆`: [u8(0xF8), 0x87] // U+8246 <cjk>
	`艉`: [u8(0xF8), 0x88] // U+8249 <cjk>
	`艅`: [u8(0xF8), 0x89] // U+8245 <cjk>
	`𦩘`: [u8(0xF8), 0x8A] // U+26A58 <cjk>
	`艋`: [u8(0xF8), 0x8B] // U+824B <cjk>
	`䑶`: [u8(0xF8), 0x8C] // U+4476 <cjk>
	`艏`: [u8(0xF8), 0x8D] // U+824F <cjk>
	`䑺`: [u8(0xF8), 0x8E] // U+447A <cjk>
	`艗`: [u8(0xF8), 0x8F] // U+8257 <cjk>
	`𦪌`: [u8(0xF8), 0x90] // U+26A8C <cjk>
	`艜`: [u8(0xF8), 0x91] // U+825C <cjk>
	`艣`: [u8(0xF8), 0x92] // U+8263 <cjk>
	`𦪷`: [u8(0xF8), 0x93] // U+26AB7 <cjk>
	`艹`: [u8(0xF8), 0x94] // U+FA5D CJK COMPATIBILITY IDEOGRAPH-FA5D
	`艹`: [u8(0xF8), 0x95] // U+FA5E CJK COMPATIBILITY IDEOGRAPH-FA5E
	`艹`: [u8(0xF8), 0x96] // U+8279 <cjk>
	`䒑`: [u8(0xF8), 0x97] // U+4491 <cjk>
	`艽`: [u8(0xF8), 0x98] // U+827D <cjk>
	`艿`: [u8(0xF8), 0x99] // U+827F <cjk>
	`芃`: [u8(0xF8), 0x9A] // U+8283 <cjk>
	`芊`: [u8(0xF8), 0x9B] // U+828A <cjk>
	`芓`: [u8(0xF8), 0x9C] // U+8293 <cjk>
	`芧`: [u8(0xF8), 0x9D] // U+82A7 <cjk>
	`芨`: [u8(0xF8), 0x9E] // U+82A8 <cjk>
	`芲`: [u8(0xF8), 0x9F] // U+82B2 <cjk>
	`芴`: [u8(0xF8), 0xA0] // U+82B4 <cjk>
	`芺`: [u8(0xF8), 0xA1] // U+82BA <cjk>
	`芼`: [u8(0xF8), 0xA2] // U+82BC <cjk>
	`苢`: [u8(0xF8), 0xA3] // U+82E2 <cjk>
	`苨`: [u8(0xF8), 0xA4] // U+82E8 <cjk>
	`苷`: [u8(0xF8), 0xA5] // U+82F7 <cjk>
	`茇`: [u8(0xF8), 0xA6] // U+8307 <cjk>
	`茈`: [u8(0xF8), 0xA7] // U+8308 <cjk>
	`茌`: [u8(0xF8), 0xA8] // U+830C <cjk>
	`荔`: [u8(0xF8), 0xA9] // U+8354 <cjk>
	`茛`: [u8(0xF8), 0xAA] // U+831B <cjk>
	`茝`: [u8(0xF8), 0xAB] // U+831D <cjk>
	`茰`: [u8(0xF8), 0xAC] // U+8330 <cjk>
	`茼`: [u8(0xF8), 0xAD] // U+833C <cjk>
	`荄`: [u8(0xF8), 0xAE] // U+8344 <cjk>
	`荗`: [u8(0xF8), 0xAF] // U+8357 <cjk>
	`䒾`: [u8(0xF8), 0xB0] // U+44BE <cjk>
	`荿`: [u8(0xF8), 0xB1] // U+837F <cjk>
	`䓔`: [u8(0xF8), 0xB2] // U+44D4 <cjk>
	`䒳`: [u8(0xF8), 0xB3] // U+44B3 <cjk>
	`莍`: [u8(0xF8), 0xB4] // U+838D <cjk>
	`莔`: [u8(0xF8), 0xB5] // U+8394 <cjk>
	`莕`: [u8(0xF8), 0xB6] // U+8395 <cjk>
	`莛`: [u8(0xF8), 0xB7] // U+839B <cjk>
	`莝`: [u8(0xF8), 0xB8] // U+839D <cjk>
	`菉`: [u8(0xF8), 0xB9] // U+83C9 <cjk>
	`菐`: [u8(0xF8), 0xBA] // U+83D0 <cjk>
	`菔`: [u8(0xF8), 0xBB] // U+83D4 <cjk>
	`菝`: [u8(0xF8), 0xBC] // U+83DD <cjk>
	`菥`: [u8(0xF8), 0xBD] // U+83E5 <cjk>
	`菹`: [u8(0xF8), 0xBE] // U+83F9 <cjk>
	`萏`: [u8(0xF8), 0xBF] // U+840F <cjk>
	`萑`: [u8(0xF8), 0xC0] // U+8411 <cjk>
	`萕`: [u8(0xF8), 0xC1] // U+8415 <cjk>
	`𦱳`: [u8(0xF8), 0xC2] // U+26C73 <cjk>
	`萗`: [u8(0xF8), 0xC3] // U+8417 <cjk>
	`萹`: [u8(0xF8), 0xC4] // U+8439 <cjk>
	`葊`: [u8(0xF8), 0xC5] // U+844A <cjk>
	`葏`: [u8(0xF8), 0xC6] // U+844F <cjk>
	`葑`: [u8(0xF8), 0xC7] // U+8451 <cjk>
	`葒`: [u8(0xF8), 0xC8] // U+8452 <cjk>
	`葙`: [u8(0xF8), 0xC9] // U+8459 <cjk>
	`葚`: [u8(0xF8), 0xCA] // U+845A <cjk>
	`葜`: [u8(0xF8), 0xCB] // U+845C <cjk>
	`𦳝`: [u8(0xF8), 0xCC] // U+26CDD <cjk>
	`葥`: [u8(0xF8), 0xCD] // U+8465 <cjk>
	`葶`: [u8(0xF8), 0xCE] // U+8476 <cjk>
	`葸`: [u8(0xF8), 0xCF] // U+8478 <cjk>
	`葼`: [u8(0xF8), 0xD0] // U+847C <cjk>
	`蒁`: [u8(0xF8), 0xD1] // U+8481 <cjk>
	`䔍`: [u8(0xF8), 0xD2] // U+450D <cjk>
	`蓜`: [u8(0xF8), 0xD3] // U+84DC <cjk>
	`蒗`: [u8(0xF8), 0xD4] // U+8497 <cjk>
	`蒦`: [u8(0xF8), 0xD5] // U+84A6 <cjk>
	`蒾`: [u8(0xF8), 0xD6] // U+84BE <cjk>
	`䔈`: [u8(0xF8), 0xD7] // U+4508 <cjk>
	`蓎`: [u8(0xF8), 0xD8] // U+84CE <cjk>
	`蓏`: [u8(0xF8), 0xD9] // U+84CF <cjk>
	`蓓`: [u8(0xF8), 0xDA] // U+84D3 <cjk>
	`𦹥`: [u8(0xF8), 0xDB] // U+26E65 <cjk>
	`蓧`: [u8(0xF8), 0xDC] // U+84E7 <cjk>
	`蓪`: [u8(0xF8), 0xDD] // U+84EA <cjk>
	`蓯`: [u8(0xF8), 0xDE] // U+84EF <cjk>
	`蓰`: [u8(0xF8), 0xDF] // U+84F0 <cjk>
	`蓱`: [u8(0xF8), 0xE0] // U+84F1 <cjk>
	`蓺`: [u8(0xF8), 0xE1] // U+84FA <cjk>
	`蓽`: [u8(0xF8), 0xE2] // U+84FD <cjk>
	`蔌`: [u8(0xF8), 0xE3] // U+850C <cjk>
	`蔛`: [u8(0xF8), 0xE4] // U+851B <cjk>
	`蔤`: [u8(0xF8), 0xE5] // U+8524 <cjk>
	`蔥`: [u8(0xF8), 0xE6] // U+8525 <cjk>
	`蔫`: [u8(0xF8), 0xE7] // U+852B <cjk>
	`蔴`: [u8(0xF8), 0xE8] // U+8534 <cjk>
	`蕏`: [u8(0xF8), 0xE9] // U+854F <cjk>
	`蕯`: [u8(0xF8), 0xEA] // U+856F <cjk>
	`䔥`: [u8(0xF8), 0xEB] // U+4525 <cjk>
	`䕃`: [u8(0xF8), 0xEC] // U+4543 <cjk>
	`蔾`: [u8(0xF8), 0xED] // U+853E <cjk>
	`蕑`: [u8(0xF8), 0xEE] // U+8551 <cjk>
	`蕓`: [u8(0xF8), 0xEF] // U+8553 <cjk>
	`蕞`: [u8(0xF8), 0xF0] // U+855E <cjk>
	`蕡`: [u8(0xF8), 0xF1] // U+8561 <cjk>
	`蕢`: [u8(0xF8), 0xF2] // U+8562 <cjk>
	`𦾔`: [u8(0xF8), 0xF3] // U+26F94 <cjk>
	`蕻`: [u8(0xF8), 0xF4] // U+857B <cjk>
	`蕽`: [u8(0xF8), 0xF5] // U+857D <cjk>
	`蕿`: [u8(0xF8), 0xF6] // U+857F <cjk>
	`薁`: [u8(0xF8), 0xF7] // U+8581 <cjk>
	`薆`: [u8(0xF8), 0xF8] // U+8586 <cjk>
	`薓`: [u8(0xF8), 0xF9] // U+8593 <cjk>
	`薝`: [u8(0xF8), 0xFA] // U+859D <cjk>
	`薟`: [u8(0xF8), 0xFB] // U+859F <cjk>
	`𦿸`: [u8(0xF8), 0xFC] // U+26FF8 <cjk>
	`𦿶`: [u8(0xF9), 0x40] // U+26FF6 <cjk>
	`𦿷`: [u8(0xF9), 0x41] // U+26FF7 <cjk>
	`薷`: [u8(0xF9), 0x42] // U+85B7 <cjk>
	`薼`: [u8(0xF9), 0x43] // U+85BC <cjk>
	`藇`: [u8(0xF9), 0x44] // U+85C7 <cjk>
	`藊`: [u8(0xF9), 0x45] // U+85CA <cjk>
	`藘`: [u8(0xF9), 0x46] // U+85D8 <cjk>
	`藙`: [u8(0xF9), 0x47] // U+85D9 <cjk>
	`藟`: [u8(0xF9), 0x48] // U+85DF <cjk>
	`藡`: [u8(0xF9), 0x49] // U+85E1 <cjk>
	`藦`: [u8(0xF9), 0x4A] // U+85E6 <cjk>
	`藶`: [u8(0xF9), 0x4B] // U+85F6 <cjk>
	`蘀`: [u8(0xF9), 0x4C] // U+8600 <cjk>
	`蘑`: [u8(0xF9), 0x4D] // U+8611 <cjk>
	`蘞`: [u8(0xF9), 0x4E] // U+861E <cjk>
	`蘡`: [u8(0xF9), 0x4F] // U+8621 <cjk>
	`蘤`: [u8(0xF9), 0x50] // U+8624 <cjk>
	`蘧`: [u8(0xF9), 0x51] // U+8627 <cjk>
	`𧄍`: [u8(0xF9), 0x52] // U+2710D <cjk>
	`蘹`: [u8(0xF9), 0x53] // U+8639 <cjk>
	`蘼`: [u8(0xF9), 0x54] // U+863C <cjk>
	`𧄹`: [u8(0xF9), 0x55] // U+27139 <cjk>
	`虀`: [u8(0xF9), 0x56] // U+8640 <cjk>
	`蘒`: [u8(0xF9), 0x57] // U+FA20 CJK COMPATIBILITY IDEOGRAPH-FA20
	`虓`: [u8(0xF9), 0x58] // U+8653 <cjk>
	`虖`: [u8(0xF9), 0x59] // U+8656 <cjk>
	`虯`: [u8(0xF9), 0x5A] // U+866F <cjk>
	`虷`: [u8(0xF9), 0x5B] // U+8677 <cjk>
	`虺`: [u8(0xF9), 0x5C] // U+867A <cjk>
	`蚇`: [u8(0xF9), 0x5D] // U+8687 <cjk>
	`蚉`: [u8(0xF9), 0x5E] // U+8689 <cjk>
	`蚍`: [u8(0xF9), 0x5F] // U+868D <cjk>
	`蚑`: [u8(0xF9), 0x60] // U+8691 <cjk>
	`蚜`: [u8(0xF9), 0x61] // U+869C <cjk>
	`蚝`: [u8(0xF9), 0x62] // U+869D <cjk>
	`蚨`: [u8(0xF9), 0x63] // U+86A8 <cjk>
	`﨡`: [u8(0xF9), 0x64] // U+FA21 CJK COMPATIBILITY IDEOGRAPH-FA21
	`蚱`: [u8(0xF9), 0x65] // U+86B1 <cjk>
	`蚳`: [u8(0xF9), 0x66] // U+86B3 <cjk>
	`蛁`: [u8(0xF9), 0x67] // U+86C1 <cjk>
	`蛃`: [u8(0xF9), 0x68] // U+86C3 <cjk>
	`蛑`: [u8(0xF9), 0x69] // U+86D1 <cjk>
	`蛕`: [u8(0xF9), 0x6A] // U+86D5 <cjk>
	`蛗`: [u8(0xF9), 0x6B] // U+86D7 <cjk>
	`蛣`: [u8(0xF9), 0x6C] // U+86E3 <cjk>
	`蛦`: [u8(0xF9), 0x6D] // U+86E6 <cjk>
	`䖸`: [u8(0xF9), 0x6E] // U+45B8 <cjk>
	`蜅`: [u8(0xF9), 0x6F] // U+8705 <cjk>
	`蜇`: [u8(0xF9), 0x70] // U+8707 <cjk>
	`蜎`: [u8(0xF9), 0x71] // U+870E <cjk>
	`蜐`: [u8(0xF9), 0x72] // U+8710 <cjk>
	`蜓`: [u8(0xF9), 0x73] // U+8713 <cjk>
	`蜙`: [u8(0xF9), 0x74] // U+8719 <cjk>
	`蜟`: [u8(0xF9), 0x75] // U+871F <cjk>
	`蜡`: [u8(0xF9), 0x76] // U+8721 <cjk>
	`蜣`: [u8(0xF9), 0x77] // U+8723 <cjk>
	`蜱`: [u8(0xF9), 0x78] // U+8731 <cjk>
	`蜺`: [u8(0xF9), 0x79] // U+873A <cjk>
	`蜾`: [u8(0xF9), 0x7A] // U+873E <cjk>
	`蝀`: [u8(0xF9), 0x7B] // U+8740 <cjk>
	`蝃`: [u8(0xF9), 0x7C] // U+8743 <cjk>
	`蝑`: [u8(0xF9), 0x7D] // U+8751 <cjk>
	`蝘`: [u8(0xF9), 0x7E] // U+8758 <cjk>
	`蝤`: [u8(0xF9), 0x80] // U+8764 <cjk>
	`蝥`: [u8(0xF9), 0x81] // U+8765 <cjk>
	`蝲`: [u8(0xF9), 0x82] // U+8772 <cjk>
	`蝼`: [u8(0xF9), 0x83] // U+877C <cjk>
	`𧏛`: [u8(0xF9), 0x84] // U+273DB <cjk>
	`𧏚`: [u8(0xF9), 0x85] // U+273DA <cjk>
	`螧`: [u8(0xF9), 0x86] // U+87A7 <cjk>
	`螉`: [u8(0xF9), 0x87] // U+8789 <cjk>
	`螋`: [u8(0xF9), 0x88] // U+878B <cjk>
	`螓`: [u8(0xF9), 0x89] // U+8793 <cjk>
	`螠`: [u8(0xF9), 0x8A] // U+87A0 <cjk>
	`𧏾`: [u8(0xF9), 0x8B] // U+273FE <cjk>
	`䗥`: [u8(0xF9), 0x8C] // U+45E5 <cjk>
	`螾`: [u8(0xF9), 0x8D] // U+87BE <cjk>
	`𧐐`: [u8(0xF9), 0x8E] // U+27410 <cjk>
	`蟁`: [u8(0xF9), 0x8F] // U+87C1 <cjk>
	`蟎`: [u8(0xF9), 0x90] // U+87CE <cjk>
	`蟵`: [u8(0xF9), 0x91] // U+87F5 <cjk>
	`蟟`: [u8(0xF9), 0x92] // U+87DF <cjk>
	`𧑉`: [u8(0xF9), 0x93] // U+27449 <cjk>
	`蟣`: [u8(0xF9), 0x94] // U+87E3 <cjk>
	`蟥`: [u8(0xF9), 0x95] // U+87E5 <cjk>
	`蟦`: [u8(0xF9), 0x96] // U+87E6 <cjk>
	`蟪`: [u8(0xF9), 0x97] // U+87EA <cjk>
	`蟫`: [u8(0xF9), 0x98] // U+87EB <cjk>
	`蟭`: [u8(0xF9), 0x99] // U+87ED <cjk>
	`蠁`: [u8(0xF9), 0x9A] // U+8801 <cjk>
	`蠃`: [u8(0xF9), 0x9B] // U+8803 <cjk>
	`蠋`: [u8(0xF9), 0x9C] // U+880B <cjk>
	`蠓`: [u8(0xF9), 0x9D] // U+8813 <cjk>
	`蠨`: [u8(0xF9), 0x9E] // U+8828 <cjk>
	`蠮`: [u8(0xF9), 0x9F] // U+882E <cjk>
	`蠲`: [u8(0xF9), 0xA0] // U+8832 <cjk>
	`蠼`: [u8(0xF9), 0xA1] // U+883C <cjk>
	`䘏`: [u8(0xF9), 0xA2] // U+460F <cjk>
	`衊`: [u8(0xF9), 0xA3] // U+884A <cjk>
	`衘`: [u8(0xF9), 0xA4] // U+8858 <cjk>
	`衟`: [u8(0xF9), 0xA5] // U+885F <cjk>
	`衤`: [u8(0xF9), 0xA6] // U+8864 <cjk>
	`𧘕`: [u8(0xF9), 0xA7] // U+27615 <cjk>
	`𧘔`: [u8(0xF9), 0xA8] // U+27614 <cjk>
	`衩`: [u8(0xF9), 0xA9] // U+8869 <cjk>
	`𧘱`: [u8(0xF9), 0xAA] // U+27631 <cjk>
	`衯`: [u8(0xF9), 0xAB] // U+886F <cjk>
	`袠`: [u8(0xF9), 0xAC] // U+88A0 <cjk>
	`袼`: [u8(0xF9), 0xAD] // U+88BC <cjk>
	`袽`: [u8(0xF9), 0xAE] // U+88BD <cjk>
	`袾`: [u8(0xF9), 0xAF] // U+88BE <cjk>
	`裀`: [u8(0xF9), 0xB0] // U+88C0 <cjk>
	`裒`: [u8(0xF9), 0xB1] // U+88D2 <cjk>
	`𧚓`: [u8(0xF9), 0xB2] // U+27693 <cjk>
	`裑`: [u8(0xF9), 0xB3] // U+88D1 <cjk>
	`裓`: [u8(0xF9), 0xB4] // U+88D3 <cjk>
	`裛`: [u8(0xF9), 0xB5] // U+88DB <cjk>
	`裰`: [u8(0xF9), 0xB6] // U+88F0 <cjk>
	`裱`: [u8(0xF9), 0xB7] // U+88F1 <cjk>
	`䙁`: [u8(0xF9), 0xB8] // U+4641 <cjk>
	`褁`: [u8(0xF9), 0xB9] // U+8901 <cjk>
	`𧜎`: [u8(0xF9), 0xBA] // U+2770E <cjk>
	`褷`: [u8(0xF9), 0xBB] // U+8937 <cjk>
	`𧜣`: [u8(0xF9), 0xBC] // U+27723 <cjk>
	`襂`: [u8(0xF9), 0xBD] // U+8942 <cjk>
	`襅`: [u8(0xF9), 0xBE] // U+8945 <cjk>
	`襉`: [u8(0xF9), 0xBF] // U+8949 <cjk>
	`𧝒`: [u8(0xF9), 0xC0] // U+27752 <cjk>
	`䙥`: [u8(0xF9), 0xC1] // U+4665 <cjk>
	`襢`: [u8(0xF9), 0xC2] // U+8962 <cjk>
	`覀`: [u8(0xF9), 0xC3] // U+8980 <cjk>
	`覉`: [u8(0xF9), 0xC4] // U+8989 <cjk>
	`覐`: [u8(0xF9), 0xC5] // U+8990 <cjk>
	`覟`: [u8(0xF9), 0xC6] // U+899F <cjk>
	`覰`: [u8(0xF9), 0xC7] // U+89B0 <cjk>
	`覷`: [u8(0xF9), 0xC8] // U+89B7 <cjk>
	`觖`: [u8(0xF9), 0xC9] // U+89D6 <cjk>
	`觘`: [u8(0xF9), 0xCA] // U+89D8 <cjk>
	`觫`: [u8(0xF9), 0xCB] // U+89EB <cjk>
	`䚡`: [u8(0xF9), 0xCC] // U+46A1 <cjk>
	`觱`: [u8(0xF9), 0xCD] // U+89F1 <cjk>
	`觳`: [u8(0xF9), 0xCE] // U+89F3 <cjk>
	`觽`: [u8(0xF9), 0xCF] // U+89FD <cjk>
	`觿`: [u8(0xF9), 0xD0] // U+89FF <cjk>
	`䚯`: [u8(0xF9), 0xD1] // U+46AF <cjk>
	`訑`: [u8(0xF9), 0xD2] // U+8A11 <cjk>
	`訔`: [u8(0xF9), 0xD3] // U+8A14 <cjk>
	`𧦅`: [u8(0xF9), 0xD4] // U+27985 <cjk>
	`訡`: [u8(0xF9), 0xD5] // U+8A21 <cjk>
	`訵`: [u8(0xF9), 0xD6] // U+8A35 <cjk>
	`訾`: [u8(0xF9), 0xD7] // U+8A3E <cjk>
	`詅`: [u8(0xF9), 0xD8] // U+8A45 <cjk>
	`詍`: [u8(0xF9), 0xD9] // U+8A4D <cjk>
	`詘`: [u8(0xF9), 0xDA] // U+8A58 <cjk>
	`誮`: [u8(0xF9), 0xDB] // U+8AAE <cjk>
	`誐`: [u8(0xF9), 0xDC] // U+8A90 <cjk>
	`誷`: [u8(0xF9), 0xDD] // U+8AB7 <cjk>
	`誾`: [u8(0xF9), 0xDE] // U+8ABE <cjk>
	`諗`: [u8(0xF9), 0xDF] // U+8AD7 <cjk>
	`諼`: [u8(0xF9), 0xE0] // U+8AFC <cjk>
	`𧪄`: [u8(0xF9), 0xE1] // U+27A84 <cjk>
	`謊`: [u8(0xF9), 0xE2] // U+8B0A <cjk>
	`謅`: [u8(0xF9), 0xE3] // U+8B05 <cjk>
	`謍`: [u8(0xF9), 0xE4] // U+8B0D <cjk>
	`謜`: [u8(0xF9), 0xE5] // U+8B1C <cjk>
	`謟`: [u8(0xF9), 0xE6] // U+8B1F <cjk>
	`謭`: [u8(0xF9), 0xE7] // U+8B2D <cjk>
	`譃`: [u8(0xF9), 0xE8] // U+8B43 <cjk>
	`䜌`: [u8(0xF9), 0xE9] // U+470C <cjk>
	`譑`: [u8(0xF9), 0xEA] // U+8B51 <cjk>
	`譞`: [u8(0xF9), 0xEB] // U+8B5E <cjk>
	`譶`: [u8(0xF9), 0xEC] // U+8B76 <cjk>
	`譿`: [u8(0xF9), 0xED] // U+8B7F <cjk>
	`讁`: [u8(0xF9), 0xEE] // U+8B81 <cjk>
	`讋`: [u8(0xF9), 0xEF] // U+8B8B <cjk>
	`讔`: [u8(0xF9), 0xF0] // U+8B94 <cjk>
	`讕`: [u8(0xF9), 0xF1] // U+8B95 <cjk>
	`讜`: [u8(0xF9), 0xF2] // U+8B9C <cjk>
	`讞`: [u8(0xF9), 0xF3] // U+8B9E <cjk>
	`谹`: [u8(0xF9), 0xF4] // U+8C39 <cjk>
	`𧮳`: [u8(0xF9), 0xF5] // U+27BB3 <cjk>
	`谽`: [u8(0xF9), 0xF6] // U+8C3D <cjk>
	`𧮾`: [u8(0xF9), 0xF7] // U+27BBE <cjk>
	`𧯇`: [u8(0xF9), 0xF8] // U+27BC7 <cjk>
	`豅`: [u8(0xF9), 0xF9] // U+8C45 <cjk>
	`豇`: [u8(0xF9), 0xFA] // U+8C47 <cjk>
	`豏`: [u8(0xF9), 0xFB] // U+8C4F <cjk>
	`豔`: [u8(0xF9), 0xFC] // U+8C54 <cjk>
	`豗`: [u8(0xFA), 0x40] // U+8C57 <cjk>
	`豩`: [u8(0xFA), 0x41] // U+8C69 <cjk>
	`豭`: [u8(0xFA), 0x42] // U+8C6D <cjk>
	`豳`: [u8(0xFA), 0x43] // U+8C73 <cjk>
	`𧲸`: [u8(0xFA), 0x44] // U+27CB8 <cjk>
	`貓`: [u8(0xFA), 0x45] // U+8C93 <cjk>
	`貒`: [u8(0xFA), 0x46] // U+8C92 <cjk>
	`貙`: [u8(0xFA), 0x47] // U+8C99 <cjk>
	`䝤`: [u8(0xFA), 0x48] // U+4764 <cjk>
	`貛`: [u8(0xFA), 0x49] // U+8C9B <cjk>
	`貤`: [u8(0xFA), 0x4A] // U+8CA4 <cjk>
	`賖`: [u8(0xFA), 0x4B] // U+8CD6 <cjk>
	`賕`: [u8(0xFA), 0x4C] // U+8CD5 <cjk>
	`賙`: [u8(0xFA), 0x4D] // U+8CD9 <cjk>
	`𧶠`: [u8(0xFA), 0x4E] // U+27DA0 <cjk>
	`賰`: [u8(0xFA), 0x4F] // U+8CF0 <cjk>
	`賱`: [u8(0xFA), 0x50] // U+8CF1 <cjk>
	`𧸐`: [u8(0xFA), 0x51] // U+27E10 <cjk>
	`贉`: [u8(0xFA), 0x52] // U+8D09 <cjk>
	`贎`: [u8(0xFA), 0x53] // U+8D0E <cjk>
	`赬`: [u8(0xFA), 0x54] // U+8D6C <cjk>
	`趄`: [u8(0xFA), 0x55] // U+8D84 <cjk>
	`趕`: [u8(0xFA), 0x56] // U+8D95 <cjk>
	`趦`: [u8(0xFA), 0x57] // U+8DA6 <cjk>
	`𧾷`: [u8(0xFA), 0x58] // U+27FB7 <cjk>
	`跆`: [u8(0xFA), 0x59] // U+8DC6 <cjk>
	`跈`: [u8(0xFA), 0x5A] // U+8DC8 <cjk>
	`跙`: [u8(0xFA), 0x5B] // U+8DD9 <cjk>
	`跬`: [u8(0xFA), 0x5C] // U+8DEC <cjk>
	`踌`: [u8(0xFA), 0x5D] // U+8E0C <cjk>
	`䟽`: [u8(0xFA), 0x5E] // U+47FD <cjk>
	`跽`: [u8(0xFA), 0x5F] // U+8DFD <cjk>
	`踆`: [u8(0xFA), 0x60] // U+8E06 <cjk>
	`𨂊`: [u8(0xFA), 0x61] // U+2808A <cjk>
	`踔`: [u8(0xFA), 0x62] // U+8E14 <cjk>
	`踖`: [u8(0xFA), 0x63] // U+8E16 <cjk>
	`踡`: [u8(0xFA), 0x64] // U+8E21 <cjk>
	`踢`: [u8(0xFA), 0x65] // U+8E22 <cjk>
	`踧`: [u8(0xFA), 0x66] // U+8E27 <cjk>
	`𨂻`: [u8(0xFA), 0x67] // U+280BB <cjk>
	`䠖`: [u8(0xFA), 0x68] // U+4816 <cjk>
	`踶`: [u8(0xFA), 0x69] // U+8E36 <cjk>
	`踹`: [u8(0xFA), 0x6A] // U+8E39 <cjk>
	`蹋`: [u8(0xFA), 0x6B] // U+8E4B <cjk>
	`蹔`: [u8(0xFA), 0x6C] // U+8E54 <cjk>
	`蹢`: [u8(0xFA), 0x6D] // U+8E62 <cjk>
	`蹬`: [u8(0xFA), 0x6E] // U+8E6C <cjk>
	`蹭`: [u8(0xFA), 0x6F] // U+8E6D <cjk>
	`蹯`: [u8(0xFA), 0x70] // U+8E6F <cjk>
	`躘`: [u8(0xFA), 0x71] // U+8E98 <cjk>
	`躞`: [u8(0xFA), 0x72] // U+8E9E <cjk>
	`躮`: [u8(0xFA), 0x73] // U+8EAE <cjk>
	`躳`: [u8(0xFA), 0x74] // U+8EB3 <cjk>
	`躵`: [u8(0xFA), 0x75] // U+8EB5 <cjk>
	`躶`: [u8(0xFA), 0x76] // U+8EB6 <cjk>
	`躻`: [u8(0xFA), 0x77] // U+8EBB <cjk>
	`𨊂`: [u8(0xFA), 0x78] // U+28282 <cjk>
	`軑`: [u8(0xFA), 0x79] // U+8ED1 <cjk>
	`軔`: [u8(0xFA), 0x7A] // U+8ED4 <cjk>
	`䡎`: [u8(0xFA), 0x7B] // U+484E <cjk>
	`軹`: [u8(0xFA), 0x7C] // U+8EF9 <cjk>
	`𨋳`: [u8(0xFA), 0x7D] // U+282F3 <cjk>
	`輀`: [u8(0xFA), 0x7E] // U+8F00 <cjk>
	`輈`: [u8(0xFA), 0x80] // U+8F08 <cjk>
	`輗`: [u8(0xFA), 0x81] // U+8F17 <cjk>
	`輫`: [u8(0xFA), 0x82] // U+8F2B <cjk>
	`轀`: [u8(0xFA), 0x83] // U+8F40 <cjk>
	`轊`: [u8(0xFA), 0x84] // U+8F4A <cjk>
	`轘`: [u8(0xFA), 0x85] // U+8F58 <cjk>
	`𨐌`: [u8(0xFA), 0x86] // U+2840C <cjk>
	`辤`: [u8(0xFA), 0x87] // U+8FA4 <cjk>
	`辴`: [u8(0xFA), 0x88] // U+8FB4 <cjk>
	`辶`: [u8(0xFA), 0x89] // U+FA66 CJK COMPATIBILITY IDEOGRAPH-FA66
	`辶`: [u8(0xFA), 0x8A] // U+8FB6 <cjk>
	`𨑕`: [u8(0xFA), 0x8B] // U+28455 <cjk>
	`迁`: [u8(0xFA), 0x8C] // U+8FC1 <cjk>
	`迆`: [u8(0xFA), 0x8D] // U+8FC6 <cjk>
	`﨤`: [u8(0xFA), 0x8E] // U+FA24 CJK COMPATIBILITY IDEOGRAPH-FA24
	`迊`: [u8(0xFA), 0x8F] // U+8FCA <cjk>
	`迍`: [u8(0xFA), 0x90] // U+8FCD <cjk>
	`迓`: [u8(0xFA), 0x91] // U+8FD3 <cjk>
	`迕`: [u8(0xFA), 0x92] // U+8FD5 <cjk>
	`迠`: [u8(0xFA), 0x93] // U+8FE0 <cjk>
	`迱`: [u8(0xFA), 0x94] // U+8FF1 <cjk>
	`迵`: [u8(0xFA), 0x95] // U+8FF5 <cjk>
	`迻`: [u8(0xFA), 0x96] // U+8FFB <cjk>
	`适`: [u8(0xFA), 0x97] // U+9002 <cjk>
	`逌`: [u8(0xFA), 0x98] // U+900C <cjk>
	`逷`: [u8(0xFA), 0x99] // U+9037 <cjk>
	`𨕫`: [u8(0xFA), 0x9A] // U+2856B <cjk>
	`遃`: [u8(0xFA), 0x9B] // U+9043 <cjk>
	`遄`: [u8(0xFA), 0x9C] // U+9044 <cjk>
	`遝`: [u8(0xFA), 0x9D] // U+905D <cjk>
	`𨗈`: [u8(0xFA), 0x9E] // U+285C8 <cjk>
	`𨗉`: [u8(0xFA), 0x9F] // U+285C9 <cjk>
	`邅`: [u8(0xFA), 0xA0] // U+9085 <cjk>
	`邌`: [u8(0xFA), 0xA1] // U+908C <cjk>
	`邐`: [u8(0xFA), 0xA2] // U+9090 <cjk>
	`阝`: [u8(0xFA), 0xA3] // U+961D <cjk>
	`邡`: [u8(0xFA), 0xA4] // U+90A1 <cjk>
	`䢵`: [u8(0xFA), 0xA5] // U+48B5 <cjk>
	`邰`: [u8(0xFA), 0xA6] // U+90B0 <cjk>
	`邶`: [u8(0xFA), 0xA7] // U+90B6 <cjk>
	`郃`: [u8(0xFA), 0xA8] // U+90C3 <cjk>
	`郈`: [u8(0xFA), 0xA9] // U+90C8 <cjk>
	`𨛗`: [u8(0xFA), 0xAA] // U+286D7 <cjk>
	`郜`: [u8(0xFA), 0xAB] // U+90DC <cjk>
	`郟`: [u8(0xFA), 0xAC] // U+90DF <cjk>
	`𨛺`: [u8(0xFA), 0xAD] // U+286FA <cjk>
	`郶`: [u8(0xFA), 0xAE] // U+90F6 <cjk>
	`郲`: [u8(0xFA), 0xAF] // U+90F2 <cjk>
	`鄀`: [u8(0xFA), 0xB0] // U+9100 <cjk>
	`郫`: [u8(0xFA), 0xB1] // U+90EB <cjk>
	`郾`: [u8(0xFA), 0xB2] // U+90FE <cjk>
	`郿`: [u8(0xFA), 0xB3] // U+90FF <cjk>
	`鄄`: [u8(0xFA), 0xB4] // U+9104 <cjk>
	`鄆`: [u8(0xFA), 0xB5] // U+9106 <cjk>
	`鄘`: [u8(0xFA), 0xB6] // U+9118 <cjk>
	`鄜`: [u8(0xFA), 0xB7] // U+911C <cjk>
	`鄞`: [u8(0xFA), 0xB8] // U+911E <cjk>
	`鄷`: [u8(0xFA), 0xB9] // U+9137 <cjk>
	`鄹`: [u8(0xFA), 0xBA] // U+9139 <cjk>
	`鄺`: [u8(0xFA), 0xBB] // U+913A <cjk>
	`酆`: [u8(0xFA), 0xBC] // U+9146 <cjk>
	`酇`: [u8(0xFA), 0xBD] // U+9147 <cjk>
	`酗`: [u8(0xFA), 0xBE] // U+9157 <cjk>
	`酙`: [u8(0xFA), 0xBF] // U+9159 <cjk>
	`酡`: [u8(0xFA), 0xC0] // U+9161 <cjk>
	`酤`: [u8(0xFA), 0xC1] // U+9164 <cjk>
	`酴`: [u8(0xFA), 0xC2] // U+9174 <cjk>
	`酹`: [u8(0xFA), 0xC3] // U+9179 <cjk>
	`醅`: [u8(0xFA), 0xC4] // U+9185 <cjk>
	`醎`: [u8(0xFA), 0xC5] // U+918E <cjk>
	`醨`: [u8(0xFA), 0xC6] // U+91A8 <cjk>
	`醮`: [u8(0xFA), 0xC7] // U+91AE <cjk>
	`醳`: [u8(0xFA), 0xC8] // U+91B3 <cjk>
	`醶`: [u8(0xFA), 0xC9] // U+91B6 <cjk>
	`釃`: [u8(0xFA), 0xCA] // U+91C3 <cjk>
	`釄`: [u8(0xFA), 0xCB] // U+91C4 <cjk>
	`釚`: [u8(0xFA), 0xCC] // U+91DA <cjk>
	`𨥉`: [u8(0xFA), 0xCD] // U+28949 <cjk>
	`𨥆`: [u8(0xFA), 0xCE] // U+28946 <cjk>
	`釬`: [u8(0xFA), 0xCF] // U+91EC <cjk>
	`釮`: [u8(0xFA), 0xD0] // U+91EE <cjk>
	`鈁`: [u8(0xFA), 0xD1] // U+9201 <cjk>
	`鈊`: [u8(0xFA), 0xD2] // U+920A <cjk>
	`鈖`: [u8(0xFA), 0xD3] // U+9216 <cjk>
	`鈗`: [u8(0xFA), 0xD4] // U+9217 <cjk>
	`𨥫`: [u8(0xFA), 0xD5] // U+2896B <cjk>
	`鈳`: [u8(0xFA), 0xD6] // U+9233 <cjk>
	`鉂`: [u8(0xFA), 0xD7] // U+9242 <cjk>
	`鉇`: [u8(0xFA), 0xD8] // U+9247 <cjk>
	`鉊`: [u8(0xFA), 0xD9] // U+924A <cjk>
	`鉎`: [u8(0xFA), 0xDA] // U+924E <cjk>
	`鉑`: [u8(0xFA), 0xDB] // U+9251 <cjk>
	`鉖`: [u8(0xFA), 0xDC] // U+9256 <cjk>
	`鉙`: [u8(0xFA), 0xDD] // U+9259 <cjk>
	`鉠`: [u8(0xFA), 0xDE] // U+9260 <cjk>
	`鉡`: [u8(0xFA), 0xDF] // U+9261 <cjk>
	`鉥`: [u8(0xFA), 0xE0] // U+9265 <cjk>
	`鉧`: [u8(0xFA), 0xE1] // U+9267 <cjk>
	`鉨`: [u8(0xFA), 0xE2] // U+9268 <cjk>
	`𨦇`: [u8(0xFA), 0xE3] // U+28987 <cjk>
	`𨦈`: [u8(0xFA), 0xE4] // U+28988 <cjk>
	`鉼`: [u8(0xFA), 0xE5] // U+927C <cjk>
	`鉽`: [u8(0xFA), 0xE6] // U+927D <cjk>
	`鉿`: [u8(0xFA), 0xE7] // U+927F <cjk>
	`銉`: [u8(0xFA), 0xE8] // U+9289 <cjk>
	`銍`: [u8(0xFA), 0xE9] // U+928D <cjk>
	`銗`: [u8(0xFA), 0xEA] // U+9297 <cjk>
	`銙`: [u8(0xFA), 0xEB] // U+9299 <cjk>
	`銟`: [u8(0xFA), 0xEC] // U+929F <cjk>
	`銧`: [u8(0xFA), 0xED] // U+92A7 <cjk>
	`銫`: [u8(0xFA), 0xEE] // U+92AB <cjk>
	`𨦺`: [u8(0xFA), 0xEF] // U+289BA <cjk>
	`𨦻`: [u8(0xFA), 0xF0] // U+289BB <cjk>
	`銲`: [u8(0xFA), 0xF1] // U+92B2 <cjk>
	`銿`: [u8(0xFA), 0xF2] // U+92BF <cjk>
	`鋀`: [u8(0xFA), 0xF3] // U+92C0 <cjk>
	`鋆`: [u8(0xFA), 0xF4] // U+92C6 <cjk>
	`鋎`: [u8(0xFA), 0xF5] // U+92CE <cjk>
	`鋐`: [u8(0xFA), 0xF6] // U+92D0 <cjk>
	`鋗`: [u8(0xFA), 0xF7] // U+92D7 <cjk>
	`鋙`: [u8(0xFA), 0xF8] // U+92D9 <cjk>
	`鋥`: [u8(0xFA), 0xF9] // U+92E5 <cjk>
	`鋧`: [u8(0xFA), 0xFA] // U+92E7 <cjk>
	`錑`: [u8(0xFA), 0xFB] // U+9311 <cjk>
	`𨨞`: [u8(0xFA), 0xFC] // U+28A1E <cjk>
	`𨨩`: [u8(0xFB), 0x40] // U+28A29 <cjk>
	`鋷`: [u8(0xFB), 0x41] // U+92F7 <cjk>
	`鋹`: [u8(0xFB), 0x42] // U+92F9 <cjk>
	`鋻`: [u8(0xFB), 0x43] // U+92FB <cjk>
	`錂`: [u8(0xFB), 0x44] // U+9302 <cjk>
	`錍`: [u8(0xFB), 0x45] // U+930D <cjk>
	`錕`: [u8(0xFB), 0x46] // U+9315 <cjk>
	`錝`: [u8(0xFB), 0x47] // U+931D <cjk>
	`錞`: [u8(0xFB), 0x48] // U+931E <cjk>
	`錧`: [u8(0xFB), 0x49] // U+9327 <cjk>
	`錩`: [u8(0xFB), 0x4A] // U+9329 <cjk>
	`𨩱`: [u8(0xFB), 0x4B] // U+28A71 <cjk>
	`𨩃`: [u8(0xFB), 0x4C] // U+28A43 <cjk>
	`鍇`: [u8(0xFB), 0x4D] // U+9347 <cjk>
	`鍑`: [u8(0xFB), 0x4E] // U+9351 <cjk>
	`鍗`: [u8(0xFB), 0x4F] // U+9357 <cjk>
	`鍚`: [u8(0xFB), 0x50] // U+935A <cjk>
	`鍫`: [u8(0xFB), 0x51] // U+936B <cjk>
	`鍱`: [u8(0xFB), 0x52] // U+9371 <cjk>
	`鍳`: [u8(0xFB), 0x53] // U+9373 <cjk>
	`鎡`: [u8(0xFB), 0x54] // U+93A1 <cjk>
	`𨪙`: [u8(0xFB), 0x55] // U+28A99 <cjk>
	`𨫍`: [u8(0xFB), 0x56] // U+28ACD <cjk>
	`鎈`: [u8(0xFB), 0x57] // U+9388 <cjk>
	`鎋`: [u8(0xFB), 0x58] // U+938B <cjk>
	`鎏`: [u8(0xFB), 0x59] // U+938F <cjk>
	`鎞`: [u8(0xFB), 0x5A] // U+939E <cjk>
	`鏵`: [u8(0xFB), 0x5B] // U+93F5 <cjk>
	`𨫤`: [u8(0xFB), 0x5C] // U+28AE4 <cjk>
	`𨫝`: [u8(0xFB), 0x5D] // U+28ADD <cjk>
	`鏱`: [u8(0xFB), 0x5E] // U+93F1 <cjk>
	`鏁`: [u8(0xFB), 0x5F] // U+93C1 <cjk>
	`鏇`: [u8(0xFB), 0x60] // U+93C7 <cjk>
	`鏜`: [u8(0xFB), 0x61] // U+93DC <cjk>
	`鏢`: [u8(0xFB), 0x62] // U+93E2 <cjk>
	`鏧`: [u8(0xFB), 0x63] // U+93E7 <cjk>
	`鐉`: [u8(0xFB), 0x64] // U+9409 <cjk>
	`鐏`: [u8(0xFB), 0x65] // U+940F <cjk>
	`鐖`: [u8(0xFB), 0x66] // U+9416 <cjk>
	`鐗`: [u8(0xFB), 0x67] // U+9417 <cjk>
	`鏻`: [u8(0xFB), 0x68] // U+93FB <cjk>
	`鐲`: [u8(0xFB), 0x69] // U+9432 <cjk>
	`鐴`: [u8(0xFB), 0x6A] // U+9434 <cjk>
	`鐻`: [u8(0xFB), 0x6B] // U+943B <cjk>
	`鑅`: [u8(0xFB), 0x6C] // U+9445 <cjk>
	`𨯁`: [u8(0xFB), 0x6D] // U+28BC1 <cjk>
	`𨯯`: [u8(0xFB), 0x6E] // U+28BEF <cjk>
	`鑭`: [u8(0xFB), 0x6F] // U+946D <cjk>
	`鑯`: [u8(0xFB), 0x70] // U+946F <cjk>
	`镸`: [u8(0xFB), 0x71] // U+9578 <cjk>
	`镹`: [u8(0xFB), 0x72] // U+9579 <cjk>
	`閆`: [u8(0xFB), 0x73] // U+9586 <cjk>
	`閌`: [u8(0xFB), 0x74] // U+958C <cjk>
	`閍`: [u8(0xFB), 0x75] // U+958D <cjk>
	`𨴐`: [u8(0xFB), 0x76] // U+28D10 <cjk>
	`閫`: [u8(0xFB), 0x77] // U+95AB <cjk>
	`閴`: [u8(0xFB), 0x78] // U+95B4 <cjk>
	`𨵱`: [u8(0xFB), 0x79] // U+28D71 <cjk>
	`闈`: [u8(0xFB), 0x7A] // U+95C8 <cjk>
	`𨷻`: [u8(0xFB), 0x7B] // U+28DFB <cjk>
	`𨸟`: [u8(0xFB), 0x7C] // U+28E1F <cjk>
	`阬`: [u8(0xFB), 0x7D] // U+962C <cjk>
	`阳`: [u8(0xFB), 0x7E] // U+9633 <cjk>
	`阴`: [u8(0xFB), 0x80] // U+9634 <cjk>
	`𨸶`: [u8(0xFB), 0x81] // U+28E36 <cjk>
	`阼`: [u8(0xFB), 0x82] // U+963C <cjk>
	`陁`: [u8(0xFB), 0x83] // U+9641 <cjk>
	`陡`: [u8(0xFB), 0x84] // U+9661 <cjk>
	`𨺉`: [u8(0xFB), 0x85] // U+28E89 <cjk>
	`隂`: [u8(0xFB), 0x86] // U+9682 <cjk>
	`𨻫`: [u8(0xFB), 0x87] // U+28EEB <cjk>
	`隚`: [u8(0xFB), 0x88] // U+969A <cjk>
	`𨼲`: [u8(0xFB), 0x89] // U+28F32 <cjk>
	`䧧`: [u8(0xFB), 0x8A] // U+49E7 <cjk>
	`隩`: [u8(0xFB), 0x8B] // U+96A9 <cjk>
	`隯`: [u8(0xFB), 0x8C] // U+96AF <cjk>
	`隳`: [u8(0xFB), 0x8D] // U+96B3 <cjk>
	`隺`: [u8(0xFB), 0x8E] // U+96BA <cjk>
	`隽`: [u8(0xFB), 0x8F] // U+96BD <cjk>
	`䧺`: [u8(0xFB), 0x90] // U+49FA <cjk>
	`𨿸`: [u8(0xFB), 0x91] // U+28FF8 <cjk>
	`雘`: [u8(0xFB), 0x92] // U+96D8 <cjk>
	`雚`: [u8(0xFB), 0x93] // U+96DA <cjk>
	`雝`: [u8(0xFB), 0x94] // U+96DD <cjk>
	`䨄`: [u8(0xFB), 0x95] // U+4A04 <cjk>
	`霔`: [u8(0xFB), 0x96] // U+9714 <cjk>
	`霣`: [u8(0xFB), 0x97] // U+9723 <cjk>
	`䨩`: [u8(0xFB), 0x98] // U+4A29 <cjk>
	`霶`: [u8(0xFB), 0x99] // U+9736 <cjk>
	`靁`: [u8(0xFB), 0x9A] // U+9741 <cjk>
	`靇`: [u8(0xFB), 0x9B] // U+9747 <cjk>
	`靕`: [u8(0xFB), 0x9C] // U+9755 <cjk>
	`靗`: [u8(0xFB), 0x9D] // U+9757 <cjk>
	`靛`: [u8(0xFB), 0x9E] // U+975B <cjk>
	`靪`: [u8(0xFB), 0x9F] // U+976A <cjk>
	`𩊠`: [u8(0xFB), 0xA0] // U+292A0 <cjk>
	`𩊱`: [u8(0xFB), 0xA1] // U+292B1 <cjk>
	`鞖`: [u8(0xFB), 0xA2] // U+9796 <cjk>
	`鞚`: [u8(0xFB), 0xA3] // U+979A <cjk>
	`鞞`: [u8(0xFB), 0xA4] // U+979E <cjk>
	`鞢`: [u8(0xFB), 0xA5] // U+97A2 <cjk>
	`鞱`: [u8(0xFB), 0xA6] // U+97B1 <cjk>
	`鞲`: [u8(0xFB), 0xA7] // U+97B2 <cjk>
	`鞾`: [u8(0xFB), 0xA8] // U+97BE <cjk>
	`韌`: [u8(0xFB), 0xA9] // U+97CC <cjk>
	`韑`: [u8(0xFB), 0xAA] // U+97D1 <cjk>
	`韔`: [u8(0xFB), 0xAB] // U+97D4 <cjk>
	`韘`: [u8(0xFB), 0xAC] // U+97D8 <cjk>
	`韙`: [u8(0xFB), 0xAD] // U+97D9 <cjk>
	`韡`: [u8(0xFB), 0xAE] // U+97E1 <cjk>
	`韱`: [u8(0xFB), 0xAF] // U+97F1 <cjk>
	`頄`: [u8(0xFB), 0xB0] // U+9804 <cjk>
	`頍`: [u8(0xFB), 0xB1] // U+980D <cjk>
	`頎`: [u8(0xFB), 0xB2] // U+980E <cjk>
	`頔`: [u8(0xFB), 0xB3] // U+9814 <cjk>
	`頖`: [u8(0xFB), 0xB4] // U+9816 <cjk>
	`䪼`: [u8(0xFB), 0xB5] // U+4ABC <cjk>
	`𩒐`: [u8(0xFB), 0xB6] // U+29490 <cjk>
	`頣`: [u8(0xFB), 0xB7] // U+9823 <cjk>
	`頲`: [u8(0xFB), 0xB8] // U+9832 <cjk>
	`頳`: [u8(0xFB), 0xB9] // U+9833 <cjk>
	`頥`: [u8(0xFB), 0xBA] // U+9825 <cjk>
	`顇`: [u8(0xFB), 0xBB] // U+9847 <cjk>
	`顦`: [u8(0xFB), 0xBC] // U+9866 <cjk>
	`颫`: [u8(0xFB), 0xBD] // U+98AB <cjk>
	`颭`: [u8(0xFB), 0xBE] // U+98AD <cjk>
	`颰`: [u8(0xFB), 0xBF] // U+98B0 <cjk>
	`𩗏`: [u8(0xFB), 0xC0] // U+295CF <cjk>
	`颷`: [u8(0xFB), 0xC1] // U+98B7 <cjk>
	`颸`: [u8(0xFB), 0xC2] // U+98B8 <cjk>
	`颻`: [u8(0xFB), 0xC3] // U+98BB <cjk>
	`颼`: [u8(0xFB), 0xC4] // U+98BC <cjk>
	`颿`: [u8(0xFB), 0xC5] // U+98BF <cjk>
	`飂`: [u8(0xFB), 0xC6] // U+98C2 <cjk>
	`飇`: [u8(0xFB), 0xC7] // U+98C7 <cjk>
	`飋`: [u8(0xFB), 0xC8] // U+98CB <cjk>
	`飠`: [u8(0xFB), 0xC9] // U+98E0 <cjk>
	`𩙿`: [u8(0xFB), 0xCA] // U+2967F <cjk>
	`飡`: [u8(0xFB), 0xCB] // U+98E1 <cjk>
	`飣`: [u8(0xFB), 0xCC] // U+98E3 <cjk>
	`飥`: [u8(0xFB), 0xCD] // U+98E5 <cjk>
	`飪`: [u8(0xFB), 0xCE] // U+98EA <cjk>
	`飰`: [u8(0xFB), 0xCF] // U+98F0 <cjk>
	`飱`: [u8(0xFB), 0xD0] // U+98F1 <cjk>
	`飳`: [u8(0xFB), 0xD1] // U+98F3 <cjk>
	`餈`: [u8(0xFB), 0xD2] // U+9908 <cjk>
	`䬻`: [u8(0xFB), 0xD3] // U+4B3B <cjk>
	`𩛰`: [u8(0xFB), 0xD4] // U+296F0 <cjk>
	`餖`: [u8(0xFB), 0xD5] // U+9916 <cjk>
	`餗`: [u8(0xFB), 0xD6] // U+9917 <cjk>
	`𩜙`: [u8(0xFB), 0xD7] // U+29719 <cjk>
	`餚`: [u8(0xFB), 0xD8] // U+991A <cjk>
	`餛`: [u8(0xFB), 0xD9] // U+991B <cjk>
	`餜`: [u8(0xFB), 0xDA] // U+991C <cjk>
	`𩝐`: [u8(0xFB), 0xDB] // U+29750 <cjk>
	`餱`: [u8(0xFB), 0xDC] // U+9931 <cjk>
	`餲`: [u8(0xFB), 0xDD] // U+9932 <cjk>
	`餳`: [u8(0xFB), 0xDE] // U+9933 <cjk>
	`餺`: [u8(0xFB), 0xDF] // U+993A <cjk>
	`餻`: [u8(0xFB), 0xE0] // U+993B <cjk>
	`餼`: [u8(0xFB), 0xE1] // U+993C <cjk>
	`饀`: [u8(0xFB), 0xE2] // U+9940 <cjk>
	`饁`: [u8(0xFB), 0xE3] // U+9941 <cjk>
	`饆`: [u8(0xFB), 0xE4] // U+9946 <cjk>
	`饍`: [u8(0xFB), 0xE5] // U+994D <cjk>
	`饎`: [u8(0xFB), 0xE6] // U+994E <cjk>
	`饜`: [u8(0xFB), 0xE7] // U+995C <cjk>
	`饟`: [u8(0xFB), 0xE8] // U+995F <cjk>
	`饠`: [u8(0xFB), 0xE9] // U+9960 <cjk>
	`馣`: [u8(0xFB), 0xEA] // U+99A3 <cjk>
	`馦`: [u8(0xFB), 0xEB] // U+99A6 <cjk>
	`馹`: [u8(0xFB), 0xEC] // U+99B9 <cjk>
	`馽`: [u8(0xFB), 0xED] // U+99BD <cjk>
	`馿`: [u8(0xFB), 0xEE] // U+99BF <cjk>
	`駃`: [u8(0xFB), 0xEF] // U+99C3 <cjk>
	`駉`: [u8(0xFB), 0xF0] // U+99C9 <cjk>
	`駔`: [u8(0xFB), 0xF1] // U+99D4 <cjk>
	`駙`: [u8(0xFB), 0xF2] // U+99D9 <cjk>
	`駞`: [u8(0xFB), 0xF3] // U+99DE <cjk>
	`𩣆`: [u8(0xFB), 0xF4] // U+298C6 <cjk>
	`駰`: [u8(0xFB), 0xF5] // U+99F0 <cjk>
	`駹`: [u8(0xFB), 0xF6] // U+99F9 <cjk>
	`駼`: [u8(0xFB), 0xF7] // U+99FC <cjk>
	`騊`: [u8(0xFB), 0xF8] // U+9A0A <cjk>
	`騑`: [u8(0xFB), 0xF9] // U+9A11 <cjk>
	`騖`: [u8(0xFB), 0xFA] // U+9A16 <cjk>
	`騚`: [u8(0xFB), 0xFB] // U+9A1A <cjk>
	`騠`: [u8(0xFB), 0xFC] // U+9A20 <cjk>
	`騱`: [u8(0xFC), 0x40] // U+9A31 <cjk>
	`騶`: [u8(0xFC), 0x41] // U+9A36 <cjk>
	`驄`: [u8(0xFC), 0x42] // U+9A44 <cjk>
	`驌`: [u8(0xFC), 0x43] // U+9A4C <cjk>
	`驘`: [u8(0xFC), 0x44] // U+9A58 <cjk>
	`䯂`: [u8(0xFC), 0x45] // U+4BC2 <cjk>
	`骯`: [u8(0xFC), 0x46] // U+9AAF <cjk>
	`䯊`: [u8(0xFC), 0x47] // U+4BCA <cjk>
	`骷`: [u8(0xFC), 0x48] // U+9AB7 <cjk>
	`䯒`: [u8(0xFC), 0x49] // U+4BD2 <cjk>
	`骹`: [u8(0xFC), 0x4A] // U+9AB9 <cjk>
	`𩩲`: [u8(0xFC), 0x4B] // U+29A72 <cjk>
	`髆`: [u8(0xFC), 0x4C] // U+9AC6 <cjk>
	`髐`: [u8(0xFC), 0x4D] // U+9AD0 <cjk>
	`髒`: [u8(0xFC), 0x4E] // U+9AD2 <cjk>
	`髕`: [u8(0xFC), 0x4F] // U+9AD5 <cjk>
	`䯨`: [u8(0xFC), 0x50] // U+4BE8 <cjk>
	`髜`: [u8(0xFC), 0x51] // U+9ADC <cjk>
	`髠`: [u8(0xFC), 0x52] // U+9AE0 <cjk>
	`髥`: [u8(0xFC), 0x53] // U+9AE5 <cjk>
	`髩`: [u8(0xFC), 0x54] // U+9AE9 <cjk>
	`鬃`: [u8(0xFC), 0x55] // U+9B03 <cjk>
	`鬌`: [u8(0xFC), 0x56] // U+9B0C <cjk>
	`鬐`: [u8(0xFC), 0x57] // U+9B10 <cjk>
	`鬒`: [u8(0xFC), 0x58] // U+9B12 <cjk>
	`鬖`: [u8(0xFC), 0x59] // U+9B16 <cjk>
	`鬜`: [u8(0xFC), 0x5A] // U+9B1C <cjk>
	`鬫`: [u8(0xFC), 0x5B] // U+9B2B <cjk>
	`鬳`: [u8(0xFC), 0x5C] // U+9B33 <cjk>
	`鬽`: [u8(0xFC), 0x5D] // U+9B3D <cjk>
	`䰠`: [u8(0xFC), 0x5E] // U+4C20 <cjk>
	`魋`: [u8(0xFC), 0x5F] // U+9B4B <cjk>
	`魣`: [u8(0xFC), 0x60] // U+9B63 <cjk>
	`魥`: [u8(0xFC), 0x61] // U+9B65 <cjk>
	`魫`: [u8(0xFC), 0x62] // U+9B6B <cjk>
	`魬`: [u8(0xFC), 0x63] // U+9B6C <cjk>
	`魳`: [u8(0xFC), 0x64] // U+9B73 <cjk>
	`魶`: [u8(0xFC), 0x65] // U+9B76 <cjk>
	`魷`: [u8(0xFC), 0x66] // U+9B77 <cjk>
	`鮦`: [u8(0xFC), 0x67] // U+9BA6 <cjk>
	`鮬`: [u8(0xFC), 0x68] // U+9BAC <cjk>
	`鮱`: [u8(0xFC), 0x69] // U+9BB1 <cjk>
	`𩷛`: [u8(0xFC), 0x6A] // U+29DDB <cjk>
	`𩸽`: [u8(0xFC), 0x6B] // U+29E3D <cjk>
	`鮲`: [u8(0xFC), 0x6C] // U+9BB2 <cjk>
	`鮸`: [u8(0xFC), 0x6D] // U+9BB8 <cjk>
	`鮾`: [u8(0xFC), 0x6E] // U+9BBE <cjk>
	`鯇`: [u8(0xFC), 0x6F] // U+9BC7 <cjk>
	`鯳`: [u8(0xFC), 0x70] // U+9BF3 <cjk>
	`鯘`: [u8(0xFC), 0x71] // U+9BD8 <cjk>
	`鯝`: [u8(0xFC), 0x72] // U+9BDD <cjk>
	`鯧`: [u8(0xFC), 0x73] // U+9BE7 <cjk>
	`鯪`: [u8(0xFC), 0x74] // U+9BEA <cjk>
	`鯫`: [u8(0xFC), 0x75] // U+9BEB <cjk>
	`鯯`: [u8(0xFC), 0x76] // U+9BEF <cjk>
	`鯮`: [u8(0xFC), 0x77] // U+9BEE <cjk>
	`𩸕`: [u8(0xFC), 0x78] // U+29E15 <cjk>
	`鯺`: [u8(0xFC), 0x79] // U+9BFA <cjk>
	`𩺊`: [u8(0xFC), 0x7A] // U+29E8A <cjk>
	`鯷`: [u8(0xFC), 0x7B] // U+9BF7 <cjk>
	`𩹉`: [u8(0xFC), 0x7C] // U+29E49 <cjk>
	`鰖`: [u8(0xFC), 0x7D] // U+9C16 <cjk>
	`鰘`: [u8(0xFC), 0x7E] // U+9C18 <cjk>
	`鰙`: [u8(0xFC), 0x80] // U+9C19 <cjk>
	`鰚`: [u8(0xFC), 0x81] // U+9C1A <cjk>
	`鰝`: [u8(0xFC), 0x82] // U+9C1D <cjk>
	`鰢`: [u8(0xFC), 0x83] // U+9C22 <cjk>
	`鰧`: [u8(0xFC), 0x84] // U+9C27 <cjk>
	`鰩`: [u8(0xFC), 0x85] // U+9C29 <cjk>
	`鰪`: [u8(0xFC), 0x86] // U+9C2A <cjk>
	`𩻄`: [u8(0xFC), 0x87] // U+29EC4 <cjk>
	`鰱`: [u8(0xFC), 0x88] // U+9C31 <cjk>
	`鰶`: [u8(0xFC), 0x89] // U+9C36 <cjk>
	`鰷`: [u8(0xFC), 0x8A] // U+9C37 <cjk>
	`鱅`: [u8(0xFC), 0x8B] // U+9C45 <cjk>
	`鱜`: [u8(0xFC), 0x8C] // U+9C5C <cjk>
	`𩻩`: [u8(0xFC), 0x8D] // U+29EE9 <cjk>
	`鱉`: [u8(0xFC), 0x8E] // U+9C49 <cjk>
	`鱊`: [u8(0xFC), 0x8F] // U+9C4A <cjk>
	`𩻛`: [u8(0xFC), 0x90] // U+29EDB <cjk>
	`鱔`: [u8(0xFC), 0x91] // U+9C54 <cjk>
	`鱘`: [u8(0xFC), 0x92] // U+9C58 <cjk>
	`鱛`: [u8(0xFC), 0x93] // U+9C5B <cjk>
	`鱝`: [u8(0xFC), 0x94] // U+9C5D <cjk>
	`鱟`: [u8(0xFC), 0x95] // U+9C5F <cjk>
	`鱩`: [u8(0xFC), 0x96] // U+9C69 <cjk>
	`鱪`: [u8(0xFC), 0x97] // U+9C6A <cjk>
	`鱫`: [u8(0xFC), 0x98] // U+9C6B <cjk>
	`鱭`: [u8(0xFC), 0x99] // U+9C6D <cjk>
	`鱮`: [u8(0xFC), 0x9A] // U+9C6E <cjk>
	`鱰`: [u8(0xFC), 0x9B] // U+9C70 <cjk>
	`鱲`: [u8(0xFC), 0x9C] // U+9C72 <cjk>
	`鱵`: [u8(0xFC), 0x9D] // U+9C75 <cjk>
	`鱺`: [u8(0xFC), 0x9E] // U+9C7A <cjk>
	`鳦`: [u8(0xFC), 0x9F] // U+9CE6 <cjk>
	`鳲`: [u8(0xFC), 0xA0] // U+9CF2 <cjk>
	`鴋`: [u8(0xFC), 0xA1] // U+9D0B <cjk>
	`鴂`: [u8(0xFC), 0xA2] // U+9D02 <cjk>
	`𩿎`: [u8(0xFC), 0xA3] // U+29FCE <cjk>
	`鴑`: [u8(0xFC), 0xA4] // U+9D11 <cjk>
	`鴗`: [u8(0xFC), 0xA5] // U+9D17 <cjk>
	`鴘`: [u8(0xFC), 0xA6] // U+9D18 <cjk>
	`𪀯`: [u8(0xFC), 0xA7] // U+2A02F <cjk>
	`䳄`: [u8(0xFC), 0xA8] // U+4CC4 <cjk>
	`𪀚`: [u8(0xFC), 0xA9] // U+2A01A <cjk>
	`鴲`: [u8(0xFC), 0xAA] // U+9D32 <cjk>
	`䳑`: [u8(0xFC), 0xAB] // U+4CD1 <cjk>
	`鵂`: [u8(0xFC), 0xAC] // U+9D42 <cjk>
	`鵊`: [u8(0xFC), 0xAD] // U+9D4A <cjk>
	`鵟`: [u8(0xFC), 0xAE] // U+9D5F <cjk>
	`鵢`: [u8(0xFC), 0xAF] // U+9D62 <cjk>
	`𪃹`: [u8(0xFC), 0xB0] // U+2A0F9 <cjk>
	`鵩`: [u8(0xFC), 0xB1] // U+9D69 <cjk>
	`鵫`: [u8(0xFC), 0xB2] // U+9D6B <cjk>
	`𪂂`: [u8(0xFC), 0xB3] // U+2A082 <cjk>
	`鵳`: [u8(0xFC), 0xB4] // U+9D73 <cjk>
	`鵶`: [u8(0xFC), 0xB5] // U+9D76 <cjk>
	`鵷`: [u8(0xFC), 0xB6] // U+9D77 <cjk>
	`鵾`: [u8(0xFC), 0xB7] // U+9D7E <cjk>
	`鶄`: [u8(0xFC), 0xB8] // U+9D84 <cjk>
	`鶍`: [u8(0xFC), 0xB9] // U+9D8D <cjk>
	`鶙`: [u8(0xFC), 0xBA] // U+9D99 <cjk>
	`鶡`: [u8(0xFC), 0xBB] // U+9DA1 <cjk>
	`鶿`: [u8(0xFC), 0xBC] // U+9DBF <cjk>
	`鶵`: [u8(0xFC), 0xBD] // U+9DB5 <cjk>
	`鶹`: [u8(0xFC), 0xBE] // U+9DB9 <cjk>
	`鶽`: [u8(0xFC), 0xBF] // U+9DBD <cjk>
	`鷃`: [u8(0xFC), 0xC0] // U+9DC3 <cjk>
	`鷇`: [u8(0xFC), 0xC1] // U+9DC7 <cjk>
	`鷉`: [u8(0xFC), 0xC2] // U+9DC9 <cjk>
	`鷖`: [u8(0xFC), 0xC3] // U+9DD6 <cjk>
	`鷚`: [u8(0xFC), 0xC4] // U+9DDA <cjk>
	`鷟`: [u8(0xFC), 0xC5] // U+9DDF <cjk>
	`鷠`: [u8(0xFC), 0xC6] // U+9DE0 <cjk>
	`鷣`: [u8(0xFC), 0xC7] // U+9DE3 <cjk>
	`鷴`: [u8(0xFC), 0xC8] // U+9DF4 <cjk>
	`䴇`: [u8(0xFC), 0xC9] // U+4D07 <cjk>
	`鸊`: [u8(0xFC), 0xCA] // U+9E0A <cjk>
	`鸂`: [u8(0xFC), 0xCB] // U+9E02 <cjk>
	`鸍`: [u8(0xFC), 0xCC] // U+9E0D <cjk>
	`鸙`: [u8(0xFC), 0xCD] // U+9E19 <cjk>
	`鸜`: [u8(0xFC), 0xCE] // U+9E1C <cjk>
	`鸝`: [u8(0xFC), 0xCF] // U+9E1D <cjk>
	`鹻`: [u8(0xFC), 0xD0] // U+9E7B <cjk>
	`𢈘`: [u8(0xFC), 0xD1] // U+22218 <cjk>
	`麀`: [u8(0xFC), 0xD2] // U+9E80 <cjk>
	`麅`: [u8(0xFC), 0xD3] // U+9E85 <cjk>
	`麛`: [u8(0xFC), 0xD4] // U+9E9B <cjk>
	`麨`: [u8(0xFC), 0xD5] // U+9EA8 <cjk>
	`𪎌`: [u8(0xFC), 0xD6] // U+2A38C <cjk>
	`麽`: [u8(0xFC), 0xD7] // U+9EBD <cjk>
	`𪐷`: [u8(0xFC), 0xD8] // U+2A437 <cjk>
	`黟`: [u8(0xFC), 0xD9] // U+9EDF <cjk>
	`黧`: [u8(0xFC), 0xDA] // U+9EE7 <cjk>
	`黮`: [u8(0xFC), 0xDB] // U+9EEE <cjk>
	`黿`: [u8(0xFC), 0xDC] // U+9EFF <cjk>
	`鼂`: [u8(0xFC), 0xDD] // U+9F02 <cjk>
	`䵷`: [u8(0xFC), 0xDE] // U+4D77 <cjk>
	`鼃`: [u8(0xFC), 0xDF] // U+9F03 <cjk>
	`鼗`: [u8(0xFC), 0xE0] // U+9F17 <cjk>
	`鼙`: [u8(0xFC), 0xE1] // U+9F19 <cjk>
	`鼯`: [u8(0xFC), 0xE2] // U+9F2F <cjk>
	`鼷`: [u8(0xFC), 0xE3] // U+9F37 <cjk>
	`鼺`: [u8(0xFC), 0xE4] // U+9F3A <cjk>
	`鼽`: [u8(0xFC), 0xE5] // U+9F3D <cjk>
	`齁`: [u8(0xFC), 0xE6] // U+9F41 <cjk>
	`齅`: [u8(0xFC), 0xE7] // U+9F45 <cjk>
	`齆`: [u8(0xFC), 0xE8] // U+9F46 <cjk>
	`齓`: [u8(0xFC), 0xE9] // U+9F53 <cjk>
	`齕`: [u8(0xFC), 0xEA] // U+9F55 <cjk>
	`齘`: [u8(0xFC), 0xEB] // U+9F58 <cjk>
	`𪗱`: [u8(0xFC), 0xEC] // U+2A5F1 <cjk>
	`齝`: [u8(0xFC), 0xED] // U+9F5D <cjk>
	`𪘂`: [u8(0xFC), 0xEE] // U+2A602 <cjk>
	`齩`: [u8(0xFC), 0xEF] // U+9F69 <cjk>
	`𪘚`: [u8(0xFC), 0xF0] // U+2A61A <cjk>
	`齭`: [u8(0xFC), 0xF1] // U+9F6D <cjk>
	`齰`: [u8(0xFC), 0xF2] // U+9F70 <cjk>
	`齵`: [u8(0xFC), 0xF3] // U+9F75 <cjk>
	`𪚲`: [u8(0xFC), 0xF4] // U+2A6B2 <cjk>
}

// UTF-8 sequence for JIS X 0213
const utf8_sequence_for_jis_x_0213 = {
	'か゚': [u8(0x82), 0xF5] // U+304B+309A
	'き゚': [u8(0x82), 0xF6] // U+304D+309A
	'く゚': [u8(0x82), 0xF7] // U+304F+309A
	'け゚': [u8(0x82), 0xF8] // U+3051+309A
	'こ゚': [u8(0x82), 0xF9] // U+3053+309A
	'カ゚': [u8(0x83), 0x97] // U+30AB+309A
	'キ゚': [u8(0x83), 0x98] // U+30AD+309A
	'ク゚': [u8(0x83), 0x99] // U+30AF+309A
	'ケ゚': [u8(0x83), 0x9A] // U+30B1+309A
	'コ゚': [u8(0x83), 0x9B] // U+30B3+309A
	'セ゚': [u8(0x83), 0x9C] // U+30BB+309A
	'ツ゚': [u8(0x83), 0x9D] // U+30C4+309A
	'ト゚': [u8(0x83), 0x9E] // U+30C8+309A
	'ㇷ゚': [u8(0x83), 0xF6] // U+31F7+309A
	'æ̀': [u8(0x86), 0x63] // U+00E6+0300
	'ɔ̀': [u8(0x86), 0x67] // U+0254+0300
	'ɔ́': [u8(0x86), 0x68] // U+0254+0301
	'ʌ̀': [u8(0x86), 0x69] // U+028C+0300
	'ʌ́': [u8(0x86), 0x6A] // U+028C+0301
	'ə̀': [u8(0x86), 0x6B] // U+0259+0300
	'ə́': [u8(0x86), 0x6C] // U+0259+0301
	'ɚ̀': [u8(0x86), 0x6D] // U+025A+0300
	'ɚ́': [u8(0x86), 0x6E] // U+025A+0301
	'˩˥': [u8(0x86), 0x85] // U+02E9+02E5
	'˥˩': [u8(0x86), 0x86] // U+02E5+02E9
}

// UTF-8 possible sequences JIS X 0213
const utf8_possible_sequences_jis_x_0213 = {
	// U+309A
	`か`: [`゚`]
	`き`: [`゚`]
	`く`: [`゚`]
	`け`: [`゚`]
	`こ`: [`゚`]
	`カ`: [`゚`]
	`キ`: [`゚`]
	`ク`: [`゚`]
	`ケ`: [`゚`]
	`コ`: [`゚`]
	`セ`: [`゚`]
	`ツ`: [`゚`]
	`ト`: [`゚`]
	`ㇷ`: [`゚`]

	// U+0300; U+0301
	`æ`: [`̀`, `́`]
	`ɔ`: [`̀`, `́`]
	`ʌ`: [`̀`, `́`]
	`ə`: [`̀`, `́`]
	`ɚ`: [`̀`, `́`]

	// U+02E5; U+02E9
	`˩`: [`˥`]
	`˥`: [`˩`]
}
module mojibake

const jis_x_0213_doublebyte_0xe9 = {
	0x40: [`\u9871`].string() // U+9871 <cjk>
	0x41: [`\u9874`].string() // U+9874 <cjk>
	0x42: [`\u9873`].string() // U+9873 <cjk>
	0x43: [`\u98AA`].string() // U+98AA <cjk>
	0x44: [`\u98AF`].string() // U+98AF <cjk>
	0x45: [`\u98B1`].string() // U+98B1 <cjk>
	0x46: [`\u98B6`].string() // U+98B6 <cjk>
	0x47: [`\u98C4`].string() // U+98C4 <cjk>
	0x48: [`\u98C3`].string() // U+98C3 <cjk>
	0x49: [`\u98C6`].string() // U+98C6 <cjk>
	0x4A: [`\u98E9`].string() // U+98E9 <cjk>
	0x4B: [`\u98EB`].string() // U+98EB <cjk>
	0x4C: [`\u9903`].string() // U+9903 <cjk>
	0x4D: [`\u9909`].string() // U+9909 <cjk>
	0x4E: [`\u9912`].string() // U+9912 <cjk>
	0x4F: [`\u9914`].string() // U+9914 <cjk>
	0x50: [`\u9918`].string() // U+9918 <cjk>
	0x51: [`\u9921`].string() // U+9921 <cjk>
	0x52: [`\u991D`].string() // U+991D <cjk>
	0x53: [`\u991E`].string() // U+991E <cjk>
	0x54: [`\u9924`].string() // U+9924 <cjk>
	0x55: [`\u9920`].string() // U+9920 <cjk>
	0x56: [`\u992C`].string() // U+992C <cjk>
	0x57: [`\u992E`].string() // U+992E <cjk>
	0x58: [`\u993D`].string() // U+993D <cjk>
	0x59: [`\u993E`].string() // U+993E <cjk>
	0x5A: [`\u9942`].string() // U+9942 <cjk>
	0x5B: [`\u9949`].string() // U+9949 <cjk>
	0x5C: [`\u9945`].string() // U+9945 <cjk>
	0x5D: [`\u9950`].string() // U+9950 <cjk>
	0x5E: [`\u994B`].string() // U+994B <cjk>
	0x5F: [`\u9951`].string() // U+9951 <cjk>
	0x60: [`\u9952`].string() // U+9952 <cjk>
	0x61: [`\u994C`].string() // U+994C <cjk>
	0x62: [`\u9955`].string() // U+9955 <cjk>
	0x63: [`\u9997`].string() // U+9997 <cjk>
	0x64: [`\u9998`].string() // U+9998 <cjk>
	0x65: [`\u99A5`].string() // U+99A5 <cjk>
	0x66: [`\u99AD`].string() // U+99AD <cjk>
	0x67: [`\u99AE`].string() // U+99AE <cjk>
	0x68: [`\u99BC`].string() // U+99BC <cjk>
	0x69: [`\u99DF`].string() // U+99DF <cjk>
	0x6A: [`\u99DB`].string() // U+99DB <cjk>
	0x6B: [`\u99DD`].string() // U+99DD <cjk>
	0x6C: [`\u99D8`].string() // U+99D8 <cjk>
	0x6D: [`\u99D1`].string() // U+99D1 <cjk>
	0x6E: [`\u99ED`].string() // U+99ED <cjk>
	0x6F: [`\u99EE`].string() // U+99EE <cjk>
	0x70: [`\u99F1`].string() // U+99F1 <cjk>
	0x71: [`\u99F2`].string() // U+99F2 <cjk>
	0x72: [`\u99FB`].string() // U+99FB <cjk>
	0x73: [`\u99F8`].string() // U+99F8 <cjk>
	0x74: [`\u9A01`].string() // U+9A01 <cjk>
	0x75: [`\u9A0F`].string() // U+9A0F <cjk>
	0x76: [`\u9A05`].string() // U+9A05 <cjk>
	0x77: [`\u99E2`].string() // U+99E2 <cjk>
	0x78: [`\u9A19`].string() // U+9A19 <cjk>
	0x79: [`\u9A2B`].string() // U+9A2B <cjk>
	0x7A: [`\u9A37`].string() // U+9A37 <cjk>
	0x7B: [`\u9A45`].string() // U+9A45 <cjk>
	0x7C: [`\u9A42`].string() // U+9A42 <cjk>
	0x7D: [`\u9A40`].string() // U+9A40 <cjk>
	0x7E: [`\u9A43`].string() // U+9A43 <cjk>
	0x80: [`\u9A3E`].string() // U+9A3E <cjk>
	0x81: [`\u9A55`].string() // U+9A55 <cjk>
	0x82: [`\u9A4D`].string() // U+9A4D <cjk>
	0x83: [`\u9A5B`].string() // U+9A5B <cjk>
	0x84: [`\u9A57`].string() // U+9A57 <cjk>
	0x85: [`\u9A5F`].string() // U+9A5F <cjk>
	0x86: [`\u9A62`].string() // U+9A62 <cjk>
	0x87: [`\u9A65`].string() // U+9A65 <cjk>
	0x88: [`\u9A64`].string() // U+9A64 <cjk>
	0x89: [`\u9A69`].string() // U+9A69 <cjk>
	0x8A: [`\u9A6B`].string() // U+9A6B <cjk>
	0x8B: [`\u9A6A`].string() // U+9A6A <cjk>
	0x8C: [`\u9AAD`].string() // U+9AAD <cjk>
	0x8D: [`\u9AB0`].string() // U+9AB0 <cjk>
	0x8E: [`\u9ABC`].string() // U+9ABC <cjk>
	0x8F: [`\u9AC0`].string() // U+9AC0 <cjk>
	0x90: [`\u9ACF`].string() // U+9ACF <cjk>
	0x91: [`\u9AD1`].string() // U+9AD1 <cjk>
	0x92: [`\u9AD3`].string() // U+9AD3 <cjk>
	0x93: [`\u9AD4`].string() // U+9AD4 <cjk>
	0x94: [`\u9ADE`].string() // U+9ADE <cjk>
	0x95: [`\u9ADF`].string() // U+9ADF <cjk>
	0x96: [`\u9AE2`].string() // U+9AE2 <cjk>
	0x97: [`\u9AE3`].string() // U+9AE3 <cjk>
	0x98: [`\u9AE6`].string() // U+9AE6 <cjk>
	0x99: [`\u9AEF`].string() // U+9AEF <cjk>
	0x9A: [`\u9AEB`].string() // U+9AEB <cjk>
	0x9B: [`\u9AEE`].string() // U+9AEE <cjk>
	0x9C: [`\u9AF4`].string() // U+9AF4 <cjk>
	0x9D: [`\u9AF1`].string() // U+9AF1 <cjk>
	0x9E: [`\u9AF7`].string() // U+9AF7 <cjk>
	0x9F: [`\u9AFB`].string() // U+9AFB <cjk>
	0xA0: [`\u9B06`].string() // U+9B06 <cjk>
	0xA1: [`\u9B18`].string() // U+9B18 <cjk>
	0xA2: [`\u9B1A`].string() // U+9B1A <cjk>
	0xA3: [`\u9B1F`].string() // U+9B1F <cjk>
	0xA4: [`\u9B22`].string() // U+9B22 <cjk>
	0xA5: [`\u9B23`].string() // U+9B23 <cjk>
	0xA6: [`\u9B25`].string() // U+9B25 <cjk>
	0xA7: [`\u9B27`].string() // U+9B27 <cjk>
	0xA8: [`\u9B28`].string() // U+9B28 <cjk>
	0xA9: [`\u9B29`].string() // U+9B29 <cjk>
	0xAA: [`\u9B2A`].string() // U+9B2A <cjk>
	0xAB: [`\u9B2E`].string() // U+9B2E <cjk>
	0xAC: [`\u9B2F`].string() // U+9B2F <cjk>
	0xAD: [`\u9B32`].string() // U+9B32 <cjk>
	0xAE: [`\u9B44`].string() // U+9B44 <cjk>
	0xAF: [`\u9B43`].string() // U+9B43 <cjk>
	0xB0: [`\u9B4F`].string() // U+9B4F <cjk>
	0xB1: [`\u9B4D`].string() // U+9B4D <cjk>
	0xB2: [`\u9B4E`].string() // U+9B4E <cjk>
	0xB3: [`\u9B51`].string() // U+9B51 <cjk>
	0xB4: [`\u9B58`].string() // U+9B58 <cjk>
	0xB5: [`\u9B74`].string() // U+9B74 <cjk>
	0xB6: [`\u9B93`].string() // U+9B93 <cjk>
	0xB7: [`\u9B83`].string() // U+9B83 <cjk>
	0xB8: [`\u9B91`].string() // U+9B91 <cjk>
	0xB9: [`\u9B96`].string() // U+9B96 <cjk>
	0xBA: [`\u9B97`].string() // U+9B97 <cjk>
	0xBB: [`\u9B9F`].string() // U+9B9F <cjk>
	0xBC: [`\u9BA0`].string() // U+9BA0 <cjk>
	0xBD: [`\u9BA8`].string() // U+9BA8 <cjk>
	0xBE: [`\u9BB4`].string() // U+9BB4 <cjk>
	0xBF: [`\u9BC0`].string() // U+9BC0 <cjk>
	0xC0: [`\u9BCA`].string() // U+9BCA <cjk>
	0xC1: [`\u9BB9`].string() // U+9BB9 <cjk>
	0xC2: [`\u9BC6`].string() // U+9BC6 <cjk>
	0xC3: [`\u9BCF`].string() // U+9BCF <cjk>
	0xC4: [`\u9BD1`].string() // U+9BD1 <cjk>
	0xC5: [`\u9BD2`].string() // U+9BD2 <cjk>
	0xC6: [`\u9BE3`].string() // U+9BE3 <cjk>
	0xC7: [`\u9BE2`].string() // U+9BE2 <cjk>
	0xC8: [`\u9BE4`].string() // U+9BE4 <cjk>
	0xC9: [`\u9BD4`].string() // U+9BD4 <cjk>
	0xCA: [`\u9BE1`].string() // U+9BE1 <cjk>
	0xCB: [`\u9C3A`].string() // U+9C3A <cjk>
	0xCC: [`\u9BF2`].string() // U+9BF2 <cjk>
	0xCD: [`\u9BF1`].string() // U+9BF1 <cjk>
	0xCE: [`\u9BF0`].string() // U+9BF0 <cjk>
	0xCF: [`\u9C15`].string() // U+9C15 <cjk>
	0xD0: [`\u9C14`].string() // U+9C14 <cjk>
	0xD1: [`\u9C09`].string() // U+9C09 <cjk>
	0xD2: [`\u9C13`].string() // U+9C13 <cjk>
	0xD3: [`\u9C0C`].string() // U+9C0C <cjk>
	0xD4: [`\u9C06`].string() // U+9C06 <cjk>
	0xD5: [`\u9C08`].string() // U+9C08 <cjk>
	0xD6: [`\u9C12`].string() // U+9C12 <cjk>
	0xD7: [`\u9C0A`].string() // U+9C0A <cjk>
	0xD8: [`\u9C04`].string() // U+9C04 <cjk>
	0xD9: [`\u9C2E`].string() // U+9C2E <cjk>
	0xDA: [`\u9C1B`].string() // U+9C1B <cjk>
	0xDB: [`\u9C25`].string() // U+9C25 <cjk>
	0xDC: [`\u9C24`].string() // U+9C24 <cjk>
	0xDD: [`\u9C21`].string() // U+9C21 <cjk>
	0xDE: [`\u9C30`].string() // U+9C30 <cjk>
	0xDF: [`\u9C47`].string() // U+9C47 <cjk>
	0xE0: [`\u9C32`].string() // U+9C32 <cjk>
	0xE1: [`\u9C46`].string() // U+9C46 <cjk>
	0xE2: [`\u9C3E`].string() // U+9C3E <cjk>
	0xE3: [`\u9C5A`].string() // U+9C5A <cjk>
	0xE4: [`\u9C60`].string() // U+9C60 <cjk>
	0xE5: [`\u9C67`].string() // U+9C67 <cjk>
	0xE6: [`\u9C76`].string() // U+9C76 <cjk>
	0xE7: [`\u9C78`].string() // U+9C78 <cjk>
	0xE8: [`\u9CE7`].string() // U+9CE7 <cjk>
	0xE9: [`\u9CEC`].string() // U+9CEC <cjk>
	0xEA: [`\u9CF0`].string() // U+9CF0 <cjk>
	0xEB: [`\u9D09`].string() // U+9D09 <cjk>
	0xEC: [`\u9D08`].string() // U+9D08 <cjk>
	0xED: [`\u9CEB`].string() // U+9CEB <cjk>
	0xEE: [`\u9D03`].string() // U+9D03 <cjk>
	0xEF: [`\u9D06`].string() // U+9D06 <cjk>
	0xF0: [`\u9D2A`].string() // U+9D2A <cjk>
	0xF1: [`\u9D26`].string() // U+9D26 <cjk>
	0xF2: [`\u9DAF`].string() // U+9DAF <cjk>
	0xF3: [`\u9D23`].string() // U+9D23 <cjk>
	0xF4: [`\u9D1F`].string() // U+9D1F <cjk>
	0xF5: [`\u9D44`].string() // U+9D44 <cjk>
	0xF6: [`\u9D15`].string() // U+9D15 <cjk>
	0xF7: [`\u9D12`].string() // U+9D12 <cjk>
	0xF8: [`\u9D41`].string() // U+9D41 <cjk>
	0xF9: [`\u9D3F`].string() // U+9D3F <cjk>
	0xFA: [`\u9D3E`].string() // U+9D3E <cjk>
	0xFB: [`\u9D46`].string() // U+9D46 <cjk>
	0xFC: [`\u9D48`].string() // U+9D48 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xe8 = {
	0x40: [`\u9319`].string() // U+9319 <cjk>
	0x41: [`\u9322`].string() // U+9322 <cjk>
	0x42: [`\u931A`].string() // U+931A <cjk>
	0x43: [`\u9323`].string() // U+9323 <cjk>
	0x44: [`\u933A`].string() // U+933A <cjk>
	0x45: [`\u9335`].string() // U+9335 <cjk>
	0x46: [`\u933B`].string() // U+933B <cjk>
	0x47: [`\u935C`].string() // U+935C <cjk>
	0x48: [`\u9360`].string() // U+9360 <cjk>
	0x49: [`\u937C`].string() // U+937C <cjk>
	0x4A: [`\u936E`].string() // U+936E <cjk>
	0x4B: [`\u9356`].string() // U+9356 <cjk>
	0x4C: [`\u93B0`].string() // U+93B0 <cjk>
	0x4D: [`\u93AC`].string() // U+93AC <cjk>
	0x4E: [`\u93AD`].string() // U+93AD <cjk>
	0x4F: [`\u9394`].string() // U+9394 <cjk>
	0x50: [`\u93B9`].string() // U+93B9 <cjk>
	0x51: [`\u93D6`].string() // U+93D6 <cjk>
	0x52: [`\u93D7`].string() // U+93D7 <cjk>
	0x53: [`\u93E8`].string() // U+93E8 <cjk>
	0x54: [`\u93E5`].string() // U+93E5 <cjk>
	0x55: [`\u93D8`].string() // U+93D8 <cjk>
	0x56: [`\u93C3`].string() // U+93C3 <cjk>
	0x57: [`\u93DD`].string() // U+93DD <cjk>
	0x58: [`\u93D0`].string() // U+93D0 <cjk>
	0x59: [`\u93C8`].string() // U+93C8 <cjk>
	0x5A: [`\u93E4`].string() // U+93E4 <cjk>
	0x5B: [`\u941A`].string() // U+941A <cjk>
	0x5C: [`\u9414`].string() // U+9414 <cjk>
	0x5D: [`\u9413`].string() // U+9413 <cjk>
	0x5E: [`\u9403`].string() // U+9403 <cjk>
	0x5F: [`\u9407`].string() // U+9407 <cjk>
	0x60: [`\u9410`].string() // U+9410 <cjk>
	0x61: [`\u9436`].string() // U+9436 <cjk>
	0x62: [`\u942B`].string() // U+942B <cjk>
	0x63: [`\u9435`].string() // U+9435 <cjk>
	0x64: [`\u9421`].string() // U+9421 <cjk>
	0x65: [`\u943A`].string() // U+943A <cjk>
	0x66: [`\u9441`].string() // U+9441 <cjk>
	0x67: [`\u9452`].string() // U+9452 <cjk>
	0x68: [`\u9444`].string() // U+9444 <cjk>
	0x69: [`\u945B`].string() // U+945B <cjk>
	0x6A: [`\u9460`].string() // U+9460 <cjk>
	0x6B: [`\u9462`].string() // U+9462 <cjk>
	0x6C: [`\u945E`].string() // U+945E <cjk>
	0x6D: [`\u946A`].string() // U+946A <cjk>
	0x6E: [`\u9229`].string() // U+9229 <cjk>
	0x6F: [`\u9470`].string() // U+9470 <cjk>
	0x70: [`\u9475`].string() // U+9475 <cjk>
	0x71: [`\u9477`].string() // U+9477 <cjk>
	0x72: [`\u947D`].string() // U+947D <cjk>
	0x73: [`\u945A`].string() // U+945A <cjk>
	0x74: [`\u947C`].string() // U+947C <cjk>
	0x75: [`\u947E`].string() // U+947E <cjk>
	0x76: [`\u9481`].string() // U+9481 <cjk>
	0x77: [`\u947F`].string() // U+947F <cjk>
	0x78: [`\u9582`].string() // U+9582 <cjk>
	0x79: [`\u9587`].string() // U+9587 <cjk>
	0x7A: [`\u958A`].string() // U+958A <cjk>
	0x7B: [`\u9594`].string() // U+9594 <cjk>
	0x7C: [`\u9596`].string() // U+9596 <cjk>
	0x7D: [`\u9598`].string() // U+9598 <cjk>
	0x7E: [`\u9599`].string() // U+9599 <cjk>
	0x80: [`\u95A0`].string() // U+95A0 <cjk>
	0x81: [`\u95A8`].string() // U+95A8 <cjk>
	0x82: [`\u95A7`].string() // U+95A7 <cjk>
	0x83: [`\u95AD`].string() // U+95AD <cjk>
	0x84: [`\u95BC`].string() // U+95BC <cjk>
	0x85: [`\u95BB`].string() // U+95BB <cjk>
	0x86: [`\u95B9`].string() // U+95B9 <cjk>
	0x87: [`\u95BE`].string() // U+95BE <cjk>
	0x88: [`\u95CA`].string() // U+95CA <cjk>
	0x89: [`\u6FF6`].string() // U+6FF6 <cjk>
	0x8A: [`\u95C3`].string() // U+95C3 <cjk>
	0x8B: [`\u95CD`].string() // U+95CD <cjk>
	0x8C: [`\u95CC`].string() // U+95CC <cjk>
	0x8D: [`\u95D5`].string() // U+95D5 <cjk>
	0x8E: [`\u95D4`].string() // U+95D4 <cjk>
	0x8F: [`\u95D6`].string() // U+95D6 <cjk>
	0x90: [`\u95DC`].string() // U+95DC <cjk>
	0x91: [`\u95E1`].string() // U+95E1 <cjk>
	0x92: [`\u95E5`].string() // U+95E5 <cjk>
	0x93: [`\u95E2`].string() // U+95E2 <cjk>
	0x94: [`\u9621`].string() // U+9621 <cjk>
	0x95: [`\u9628`].string() // U+9628 <cjk>
	0x96: [`\u962E`].string() // U+962E <cjk>
	0x97: [`\u962F`].string() // U+962F <cjk>
	0x98: [`\u9642`].string() // U+9642 <cjk>
	0x99: [`\u964C`].string() // U+964C <cjk>
	0x9A: [`\u964F`].string() // U+964F <cjk>
	0x9B: [`\u964B`].string() // U+964B <cjk>
	0x9C: [`\u9677`].string() // U+9677 <cjk>
	0x9D: [`\u965C`].string() // U+965C <cjk>
	0x9E: [`\u965E`].string() // U+965E <cjk>
	0x9F: [`\u965D`].string() // U+965D <cjk>
	0xA0: [`\u965F`].string() // U+965F <cjk>
	0xA1: [`\u9666`].string() // U+9666 <cjk>
	0xA2: [`\u9672`].string() // U+9672 <cjk>
	0xA3: [`\u966C`].string() // U+966C <cjk>
	0xA4: [`\u968D`].string() // U+968D <cjk>
	0xA5: [`\u9698`].string() // U+9698 <cjk>
	0xA6: [`\u9695`].string() // U+9695 <cjk>
	0xA7: [`\u9697`].string() // U+9697 <cjk>
	0xA8: [`\u96AA`].string() // U+96AA <cjk>
	0xA9: [`\u96A7`].string() // U+96A7 <cjk>
	0xAA: [`\u96B1`].string() // U+96B1 <cjk>
	0xAB: [`\u96B2`].string() // U+96B2 <cjk>
	0xAC: [`\u96B0`].string() // U+96B0 <cjk>
	0xAD: [`\u96B4`].string() // U+96B4 <cjk>
	0xAE: [`\u96B6`].string() // U+96B6 <cjk>
	0xAF: [`\u96B8`].string() // U+96B8 <cjk>
	0xB0: [`\u96B9`].string() // U+96B9 <cjk>
	0xB1: [`\u96CE`].string() // U+96CE <cjk>
	0xB2: [`\u96CB`].string() // U+96CB <cjk>
	0xB3: [`\u96C9`].string() // U+96C9 <cjk>
	0xB4: [`\u96CD`].string() // U+96CD <cjk>
	0xB5: [`\u894D`].string() // U+894D <cjk>
	0xB6: [`\u96DC`].string() // U+96DC <cjk>
	0xB7: [`\u970D`].string() // U+970D <cjk>
	0xB8: [`\u96D5`].string() // U+96D5 <cjk>
	0xB9: [`\u96F9`].string() // U+96F9 <cjk>
	0xBA: [`\u9704`].string() // U+9704 <cjk>
	0xBB: [`\u9706`].string() // U+9706 <cjk>
	0xBC: [`\u9708`].string() // U+9708 <cjk>
	0xBD: [`\u9713`].string() // U+9713 <cjk>
	0xBE: [`\u970E`].string() // U+970E <cjk>
	0xBF: [`\u9711`].string() // U+9711 <cjk>
	0xC0: [`\u970F`].string() // U+970F <cjk>
	0xC1: [`\u9716`].string() // U+9716 <cjk>
	0xC2: [`\u9719`].string() // U+9719 <cjk>
	0xC3: [`\u9724`].string() // U+9724 <cjk>
	0xC4: [`\u972A`].string() // U+972A <cjk>
	0xC5: [`\u9730`].string() // U+9730 <cjk>
	0xC6: [`\u9739`].string() // U+9739 <cjk>
	0xC7: [`\u973D`].string() // U+973D <cjk>
	0xC8: [`\u973E`].string() // U+973E <cjk>
	0xC9: [`\u9744`].string() // U+9744 <cjk>
	0xCA: [`\u9746`].string() // U+9746 <cjk>
	0xCB: [`\u9748`].string() // U+9748 <cjk>
	0xCC: [`\u9742`].string() // U+9742 <cjk>
	0xCD: [`\u9749`].string() // U+9749 <cjk>
	0xCE: [`\u975C`].string() // U+975C <cjk>
	0xCF: [`\u9760`].string() // U+9760 <cjk>
	0xD0: [`\u9764`].string() // U+9764 <cjk>
	0xD1: [`\u9766`].string() // U+9766 <cjk>
	0xD2: [`\u9768`].string() // U+9768 <cjk>
	0xD3: [`\u52D2`].string() // U+52D2 <cjk>
	0xD4: [`\u976B`].string() // U+976B <cjk>
	0xD5: [`\u9771`].string() // U+9771 <cjk>
	0xD6: [`\u9779`].string() // U+9779 <cjk>
	0xD7: [`\u9785`].string() // U+9785 <cjk>
	0xD8: [`\u977C`].string() // U+977C <cjk>
	0xD9: [`\u9781`].string() // U+9781 <cjk>
	0xDA: [`\u977A`].string() // U+977A <cjk>
	0xDB: [`\u9786`].string() // U+9786 <cjk>
	0xDC: [`\u978B`].string() // U+978B <cjk>
	0xDD: [`\u978F`].string() // U+978F <cjk>
	0xDE: [`\u9790`].string() // U+9790 <cjk>
	0xDF: [`\u979C`].string() // U+979C <cjk>
	0xE0: [`\u97A8`].string() // U+97A8 <cjk>
	0xE1: [`\u97A6`].string() // U+97A6 <cjk>
	0xE2: [`\u97A3`].string() // U+97A3 <cjk>
	0xE3: [`\u97B3`].string() // U+97B3 <cjk>
	0xE4: [`\u97B4`].string() // U+97B4 <cjk>
	0xE5: [`\u97C3`].string() // U+97C3 <cjk>
	0xE6: [`\u97C6`].string() // U+97C6 <cjk>
	0xE7: [`\u97C8`].string() // U+97C8 <cjk>
	0xE8: [`\u97CB`].string() // U+97CB <cjk>
	0xE9: [`\u97DC`].string() // U+97DC <cjk>
	0xEA: [`\u97ED`].string() // U+97ED <cjk>
	0xEB: [`\u9F4F`].string() // U+9F4F <cjk>
	0xEC: [`\u97F2`].string() // U+97F2 <cjk>
	0xED: [`\u7ADF`].string() // U+7ADF <cjk>
	0xEE: [`\u97F6`].string() // U+97F6 <cjk>
	0xEF: [`\u97F5`].string() // U+97F5 <cjk>
	0xF0: [`\u980F`].string() // U+980F <cjk>
	0xF1: [`\u980C`].string() // U+980C <cjk>
	0xF2: [`\u9838`].string() // U+9838 <cjk>
	0xF3: [`\u9824`].string() // U+9824 <cjk>
	0xF4: [`\u9821`].string() // U+9821 <cjk>
	0xF5: [`\u9837`].string() // U+9837 <cjk>
	0xF6: [`\u983D`].string() // U+983D <cjk>
	0xF7: [`\u9846`].string() // U+9846 <cjk>
	0xF8: [`\u984F`].string() // U+984F <cjk>
	0xF9: [`\u984B`].string() // U+984B <cjk>
	0xFA: [`\u986B`].string() // U+986B <cjk>
	0xFB: [`\u986F`].string() // U+986F <cjk>
	0xFC: [`\u9870`].string() // U+9870 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0xf9 = {
	0x40: utf32_to_str(0x26FF6) // U+26FF6 <cjk>
	0x41: utf32_to_str(0x26FF7) // U+26FF7 <cjk>
	0x42: [`\u85B7`].string() // U+85B7 <cjk>
	0x43: [`\u85BC`].string() // U+85BC <cjk>
	0x44: [`\u85C7`].string() // U+85C7 <cjk>
	0x45: [`\u85CA`].string() // U+85CA <cjk>
	0x46: [`\u85D8`].string() // U+85D8 <cjk>
	0x47: [`\u85D9`].string() // U+85D9 <cjk>
	0x48: [`\u85DF`].string() // U+85DF <cjk>
	0x49: [`\u85E1`].string() // U+85E1 <cjk>
	0x4A: [`\u85E6`].string() // U+85E6 <cjk>
	0x4B: [`\u85F6`].string() // U+85F6 <cjk>
	0x4C: [`\u8600`].string() // U+8600 <cjk>
	0x4D: [`\u8611`].string() // U+8611 <cjk>
	0x4E: [`\u861E`].string() // U+861E <cjk>
	0x4F: [`\u8621`].string() // U+8621 <cjk>
	0x50: [`\u8624`].string() // U+8624 <cjk>
	0x51: [`\u8627`].string() // U+8627 <cjk>
	0x52: utf32_to_str(0x2710D) // U+2710D <cjk>
	0x53: [`\u8639`].string() // U+8639 <cjk>
	0x54: [`\u863C`].string() // U+863C <cjk>
	0x55: utf32_to_str(0x27139) // U+27139 <cjk>
	0x56: [`\u8640`].string() // U+8640 <cjk>
	0x57: [`\uFA20`].string() // U+FA20 CJK COMPATIBILITY IDEOGRAPH-FA20
	0x58: [`\u8653`].string() // U+8653 <cjk>
	0x59: [`\u8656`].string() // U+8656 <cjk>
	0x5A: [`\u866F`].string() // U+866F <cjk>
	0x5B: [`\u8677`].string() // U+8677 <cjk>
	0x5C: [`\u867A`].string() // U+867A <cjk>
	0x5D: [`\u8687`].string() // U+8687 <cjk>
	0x5E: [`\u8689`].string() // U+8689 <cjk>
	0x5F: [`\u868D`].string() // U+868D <cjk>
	0x60: [`\u8691`].string() // U+8691 <cjk>
	0x61: [`\u869C`].string() // U+869C <cjk>
	0x62: [`\u869D`].string() // U+869D <cjk>
	0x63: [`\u86A8`].string() // U+86A8 <cjk>
	0x64: [`\uFA21`].string() // U+FA21 CJK COMPATIBILITY IDEOGRAPH-FA21
	0x65: [`\u86B1`].string() // U+86B1 <cjk>
	0x66: [`\u86B3`].string() // U+86B3 <cjk>
	0x67: [`\u86C1`].string() // U+86C1 <cjk>
	0x68: [`\u86C3`].string() // U+86C3 <cjk>
	0x69: [`\u86D1`].string() // U+86D1 <cjk>
	0x6A: [`\u86D5`].string() // U+86D5 <cjk>
	0x6B: [`\u86D7`].string() // U+86D7 <cjk>
	0x6C: [`\u86E3`].string() // U+86E3 <cjk>
	0x6D: [`\u86E6`].string() // U+86E6 <cjk>
	0x6E: [`\u45B8`].string() // U+45B8 <cjk>
	0x6F: [`\u8705`].string() // U+8705 <cjk>
	0x70: [`\u8707`].string() // U+8707 <cjk>
	0x71: [`\u870E`].string() // U+870E <cjk>
	0x72: [`\u8710`].string() // U+8710 <cjk>
	0x73: [`\u8713`].string() // U+8713 <cjk>
	0x74: [`\u8719`].string() // U+8719 <cjk>
	0x75: [`\u871F`].string() // U+871F <cjk>
	0x76: [`\u8721`].string() // U+8721 <cjk>
	0x77: [`\u8723`].string() // U+8723 <cjk>
	0x78: [`\u8731`].string() // U+8731 <cjk>
	0x79: [`\u873A`].string() // U+873A <cjk>
	0x7A: [`\u873E`].string() // U+873E <cjk>
	0x7B: [`\u8740`].string() // U+8740 <cjk>
	0x7C: [`\u8743`].string() // U+8743 <cjk>
	0x7D: [`\u8751`].string() // U+8751 <cjk>
	0x7E: [`\u8758`].string() // U+8758 <cjk>
	0x80: [`\u8764`].string() // U+8764 <cjk>
	0x81: [`\u8765`].string() // U+8765 <cjk>
	0x82: [`\u8772`].string() // U+8772 <cjk>
	0x83: [`\u877C`].string() // U+877C <cjk>
	0x84: utf32_to_str(0x273DB) // U+273DB <cjk>
	0x85: utf32_to_str(0x273DA) // U+273DA <cjk>
	0x86: [`\u87A7`].string() // U+87A7 <cjk>
	0x87: [`\u8789`].string() // U+8789 <cjk>
	0x88: [`\u878B`].string() // U+878B <cjk>
	0x89: [`\u8793`].string() // U+8793 <cjk>
	0x8A: [`\u87A0`].string() // U+87A0 <cjk>
	0x8B: utf32_to_str(0x273FE) // U+273FE <cjk>
	0x8C: [`\u45E5`].string() // U+45E5 <cjk>
	0x8D: [`\u87BE`].string() // U+87BE <cjk>
	0x8E: utf32_to_str(0x27410) // U+27410 <cjk>
	0x8F: [`\u87C1`].string() // U+87C1 <cjk>
	0x90: [`\u87CE`].string() // U+87CE <cjk>
	0x91: [`\u87F5`].string() // U+87F5 <cjk>
	0x92: [`\u87DF`].string() // U+87DF <cjk>
	0x93: utf32_to_str(0x27449) // U+27449 <cjk>
	0x94: [`\u87E3`].string() // U+87E3 <cjk>
	0x95: [`\u87E5`].string() // U+87E5 <cjk>
	0x96: [`\u87E6`].string() // U+87E6 <cjk>
	0x97: [`\u87EA`].string() // U+87EA <cjk>
	0x98: [`\u87EB`].string() // U+87EB <cjk>
	0x99: [`\u87ED`].string() // U+87ED <cjk>
	0x9A: [`\u8801`].string() // U+8801 <cjk>
	0x9B: [`\u8803`].string() // U+8803 <cjk>
	0x9C: [`\u880B`].string() // U+880B <cjk>
	0x9D: [`\u8813`].string() // U+8813 <cjk>
	0x9E: [`\u8828`].string() // U+8828 <cjk>
	0x9F: [`\u882E`].string() // U+882E <cjk>
	0xA0: [`\u8832`].string() // U+8832 <cjk>
	0xA1: [`\u883C`].string() // U+883C <cjk>
	0xA2: [`\u460F`].string() // U+460F <cjk>
	0xA3: [`\u884A`].string() // U+884A <cjk>
	0xA4: [`\u8858`].string() // U+8858 <cjk>
	0xA5: [`\u885F`].string() // U+885F <cjk>
	0xA6: [`\u8864`].string() // U+8864 <cjk>
	0xA7: utf32_to_str(0x27615) // U+27615 <cjk>
	0xA8: utf32_to_str(0x27614) // U+27614 <cjk>
	0xA9: [`\u8869`].string() // U+8869 <cjk>
	0xAA: utf32_to_str(0x27631) // U+27631 <cjk>
	0xAB: [`\u886F`].string() // U+886F <cjk>
	0xAC: [`\u88A0`].string() // U+88A0 <cjk>
	0xAD: [`\u88BC`].string() // U+88BC <cjk>
	0xAE: [`\u88BD`].string() // U+88BD <cjk>
	0xAF: [`\u88BE`].string() // U+88BE <cjk>
	0xB0: [`\u88C0`].string() // U+88C0 <cjk>
	0xB1: [`\u88D2`].string() // U+88D2 <cjk>
	0xB2: utf32_to_str(0x27693) // U+27693 <cjk>
	0xB3: [`\u88D1`].string() // U+88D1 <cjk>
	0xB4: [`\u88D3`].string() // U+88D3 <cjk>
	0xB5: [`\u88DB`].string() // U+88DB <cjk>
	0xB6: [`\u88F0`].string() // U+88F0 <cjk>
	0xB7: [`\u88F1`].string() // U+88F1 <cjk>
	0xB8: [`\u4641`].string() // U+4641 <cjk>
	0xB9: [`\u8901`].string() // U+8901 <cjk>
	0xBA: utf32_to_str(0x2770E) // U+2770E <cjk>
	0xBB: [`\u8937`].string() // U+8937 <cjk>
	0xBC: utf32_to_str(0x27723) // U+27723 <cjk>
	0xBD: [`\u8942`].string() // U+8942 <cjk>
	0xBE: [`\u8945`].string() // U+8945 <cjk>
	0xBF: [`\u8949`].string() // U+8949 <cjk>
	0xC0: utf32_to_str(0x27752) // U+27752 <cjk>
	0xC1: [`\u4665`].string() // U+4665 <cjk>
	0xC2: [`\u8962`].string() // U+8962 <cjk>
	0xC3: [`\u8980`].string() // U+8980 <cjk>
	0xC4: [`\u8989`].string() // U+8989 <cjk>
	0xC5: [`\u8990`].string() // U+8990 <cjk>
	0xC6: [`\u899F`].string() // U+899F <cjk>
	0xC7: [`\u89B0`].string() // U+89B0 <cjk>
	0xC8: [`\u89B7`].string() // U+89B7 <cjk>
	0xC9: [`\u89D6`].string() // U+89D6 <cjk>
	0xCA: [`\u89D8`].string() // U+89D8 <cjk>
	0xCB: [`\u89EB`].string() // U+89EB <cjk>
	0xCC: [`\u46A1`].string() // U+46A1 <cjk>
	0xCD: [`\u89F1`].string() // U+89F1 <cjk>
	0xCE: [`\u89F3`].string() // U+89F3 <cjk>
	0xCF: [`\u89FD`].string() // U+89FD <cjk>
	0xD0: [`\u89FF`].string() // U+89FF <cjk>
	0xD1: [`\u46AF`].string() // U+46AF <cjk>
	0xD2: [`\u8A11`].string() // U+8A11 <cjk>
	0xD3: [`\u8A14`].string() // U+8A14 <cjk>
	0xD4: utf32_to_str(0x27985) // U+27985 <cjk>
	0xD5: [`\u8A21`].string() // U+8A21 <cjk>
	0xD6: [`\u8A35`].string() // U+8A35 <cjk>
	0xD7: [`\u8A3E`].string() // U+8A3E <cjk>
	0xD8: [`\u8A45`].string() // U+8A45 <cjk>
	0xD9: [`\u8A4D`].string() // U+8A4D <cjk>
	0xDA: [`\u8A58`].string() // U+8A58 <cjk>
	0xDB: [`\u8AAE`].string() // U+8AAE <cjk>
	0xDC: [`\u8A90`].string() // U+8A90 <cjk>
	0xDD: [`\u8AB7`].string() // U+8AB7 <cjk>
	0xDE: [`\u8ABE`].string() // U+8ABE <cjk>
	0xDF: [`\u8AD7`].string() // U+8AD7 <cjk>
	0xE0: [`\u8AFC`].string() // U+8AFC <cjk>
	0xE1: utf32_to_str(0x27A84) // U+27A84 <cjk>
	0xE2: [`\u8B0A`].string() // U+8B0A <cjk>
	0xE3: [`\u8B05`].string() // U+8B05 <cjk>
	0xE4: [`\u8B0D`].string() // U+8B0D <cjk>
	0xE5: [`\u8B1C`].string() // U+8B1C <cjk>
	0xE6: [`\u8B1F`].string() // U+8B1F <cjk>
	0xE7: [`\u8B2D`].string() // U+8B2D <cjk>
	0xE8: [`\u8B43`].string() // U+8B43 <cjk>
	0xE9: [`\u470C`].string() // U+470C <cjk>
	0xEA: [`\u8B51`].string() // U+8B51 <cjk>
	0xEB: [`\u8B5E`].string() // U+8B5E <cjk>
	0xEC: [`\u8B76`].string() // U+8B76 <cjk>
	0xED: [`\u8B7F`].string() // U+8B7F <cjk>
	0xEE: [`\u8B81`].string() // U+8B81 <cjk>
	0xEF: [`\u8B8B`].string() // U+8B8B <cjk>
	0xF0: [`\u8B94`].string() // U+8B94 <cjk>
	0xF1: [`\u8B95`].string() // U+8B95 <cjk>
	0xF2: [`\u8B9C`].string() // U+8B9C <cjk>
	0xF3: [`\u8B9E`].string() // U+8B9E <cjk>
	0xF4: [`\u8C39`].string() // U+8C39 <cjk>
	0xF5: utf32_to_str(0x27BB3) // U+27BB3 <cjk>
	0xF6: [`\u8C3D`].string() // U+8C3D <cjk>
	0xF7: utf32_to_str(0x27BBE) // U+27BBE <cjk>
	0xF8: utf32_to_str(0x27BC7) // U+27BC7 <cjk>
	0xF9: [`\u8C45`].string() // U+8C45 <cjk>
	0xFA: [`\u8C47`].string() // U+8C47 <cjk>
	0xFB: [`\u8C4F`].string() // U+8C4F <cjk>
	0xFC: [`\u8C54`].string() // U+8C54 <cjk>
}

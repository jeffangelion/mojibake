module mojibake

const jis_x_0213_doublebyte_0xf8 = {
	0x40: [`\u7FF2`].string() // U+7FF2 <cjk>
	0x41: [`\u8002`].string() // U+8002 <cjk>
	0x42: [`\u800A`].string() // U+800A <cjk>
	0x43: [`\u8008`].string() // U+8008 <cjk>
	0x44: [`\u800E`].string() // U+800E <cjk>
	0x45: [`\u8011`].string() // U+8011 <cjk>
	0x46: [`\u8016`].string() // U+8016 <cjk>
	0x47: [`\u8024`].string() // U+8024 <cjk>
	0x48: [`\u802C`].string() // U+802C <cjk>
	0x49: [`\u8030`].string() // U+8030 <cjk>
	0x4A: [`\u8043`].string() // U+8043 <cjk>
	0x4B: [`\u8066`].string() // U+8066 <cjk>
	0x4C: [`\u8071`].string() // U+8071 <cjk>
	0x4D: [`\u8075`].string() // U+8075 <cjk>
	0x4E: [`\u807B`].string() // U+807B <cjk>
	0x4F: [`\u8099`].string() // U+8099 <cjk>
	0x50: [`\u809C`].string() // U+809C <cjk>
	0x51: [`\u80A4`].string() // U+80A4 <cjk>
	0x52: [`\u80A7`].string() // U+80A7 <cjk>
	0x53: [`\u80B8`].string() // U+80B8 <cjk>
	0x54: utf32_to_str(0x2667E) // U+2667E <cjk>
	0x55: [`\u80C5`].string() // U+80C5 <cjk>
	0x56: [`\u80D5`].string() // U+80D5 <cjk>
	0x57: [`\u80D8`].string() // U+80D8 <cjk>
	0x58: [`\u80E6`].string() // U+80E6 <cjk>
	0x59: utf32_to_str(0x266B0) // U+266B0 <cjk>
	0x5A: [`\u810D`].string() // U+810D <cjk>
	0x5B: [`\u80F5`].string() // U+80F5 <cjk>
	0x5C: [`\u80FB`].string() // U+80FB <cjk>
	0x5D: [`\u43EE`].string() // U+43EE <cjk>
	0x5E: [`\u8135`].string() // U+8135 <cjk>
	0x5F: [`\u8116`].string() // U+8116 <cjk>
	0x60: [`\u811E`].string() // U+811E <cjk>
	0x61: [`\u43F0`].string() // U+43F0 <cjk>
	0x62: [`\u8124`].string() // U+8124 <cjk>
	0x63: [`\u8127`].string() // U+8127 <cjk>
	0x64: [`\u812C`].string() // U+812C <cjk>
	0x65: utf32_to_str(0x2671D) // U+2671D <cjk>
	0x66: [`\u813D`].string() // U+813D <cjk>
	0x67: [`\u4408`].string() // U+4408 <cjk>
	0x68: [`\u8169`].string() // U+8169 <cjk>
	0x69: [`\u4417`].string() // U+4417 <cjk>
	0x6A: [`\u8181`].string() // U+8181 <cjk>
	0x6B: [`\u441C`].string() // U+441C <cjk>
	0x6C: [`\u8184`].string() // U+8184 <cjk>
	0x6D: [`\u8185`].string() // U+8185 <cjk>
	0x6E: [`\u4422`].string() // U+4422 <cjk>
	0x6F: [`\u8198`].string() // U+8198 <cjk>
	0x70: [`\u81B2`].string() // U+81B2 <cjk>
	0x71: [`\u81C1`].string() // U+81C1 <cjk>
	0x72: [`\u81C3`].string() // U+81C3 <cjk>
	0x73: [`\u81D6`].string() // U+81D6 <cjk>
	0x74: [`\u81DB`].string() // U+81DB <cjk>
	0x75: utf32_to_str(0x268DD) // U+268DD <cjk>
	0x76: [`\u81E4`].string() // U+81E4 <cjk>
	0x77: utf32_to_str(0x268EA) // U+268EA <cjk>
	0x78: [`\u81EC`].string() // U+81EC <cjk>
	0x79: utf32_to_str(0x26951) // U+26951 <cjk>
	0x7A: [`\u81FD`].string() // U+81FD <cjk>
	0x7B: [`\u81FF`].string() // U+81FF <cjk>
	0x7C: utf32_to_str(0x2696F) // U+2696F <cjk>
	0x7D: [`\u8204`].string() // U+8204 <cjk>
	0x7E: utf32_to_str(0x269DD) // U+269DD <cjk>
	0x80: [`\u8219`].string() // U+8219 <cjk>
	0x81: [`\u8221`].string() // U+8221 <cjk>
	0x82: [`\u8222`].string() // U+8222 <cjk>
	0x83: utf32_to_str(0x26A1E) // U+26A1E <cjk>
	0x84: [`\u8232`].string() // U+8232 <cjk>
	0x85: [`\u8234`].string() // U+8234 <cjk>
	0x86: [`\u823C`].string() // U+823C <cjk>
	0x87: [`\u8246`].string() // U+8246 <cjk>
	0x88: [`\u8249`].string() // U+8249 <cjk>
	0x89: [`\u8245`].string() // U+8245 <cjk>
	0x8A: utf32_to_str(0x26A58) // U+26A58 <cjk>
	0x8B: [`\u824B`].string() // U+824B <cjk>
	0x8C: [`\u4476`].string() // U+4476 <cjk>
	0x8D: [`\u824F`].string() // U+824F <cjk>
	0x8E: [`\u447A`].string() // U+447A <cjk>
	0x8F: [`\u8257`].string() // U+8257 <cjk>
	0x90: utf32_to_str(0x26A8C) // U+26A8C <cjk>
	0x91: [`\u825C`].string() // U+825C <cjk>
	0x92: [`\u8263`].string() // U+8263 <cjk>
	0x93: utf32_to_str(0x26AB7) // U+26AB7 <cjk>
	0x94: [`\uFA5D`].string() // U+FA5D CJK COMPATIBILITY IDEOGRAPH-FA5D
	0x95: [`\uFA5E`].string() // U+FA5E CJK COMPATIBILITY IDEOGRAPH-FA5E
	0x96: [`\u8279`].string() // U+8279 <cjk>
	0x97: [`\u4491`].string() // U+4491 <cjk>
	0x98: [`\u827D`].string() // U+827D <cjk>
	0x99: [`\u827F`].string() // U+827F <cjk>
	0x9A: [`\u8283`].string() // U+8283 <cjk>
	0x9B: [`\u828A`].string() // U+828A <cjk>
	0x9C: [`\u8293`].string() // U+8293 <cjk>
	0x9D: [`\u82A7`].string() // U+82A7 <cjk>
	0x9E: [`\u82A8`].string() // U+82A8 <cjk>
	0x9F: [`\u82B2`].string() // U+82B2 <cjk>
	0xA0: [`\u82B4`].string() // U+82B4 <cjk>
	0xA1: [`\u82BA`].string() // U+82BA <cjk>
	0xA2: [`\u82BC`].string() // U+82BC <cjk>
	0xA3: [`\u82E2`].string() // U+82E2 <cjk>
	0xA4: [`\u82E8`].string() // U+82E8 <cjk>
	0xA5: [`\u82F7`].string() // U+82F7 <cjk>
	0xA6: [`\u8307`].string() // U+8307 <cjk>
	0xA7: [`\u8308`].string() // U+8308 <cjk>
	0xA8: [`\u830C`].string() // U+830C <cjk>
	0xA9: [`\u8354`].string() // U+8354 <cjk>
	0xAA: [`\u831B`].string() // U+831B <cjk>
	0xAB: [`\u831D`].string() // U+831D <cjk>
	0xAC: [`\u8330`].string() // U+8330 <cjk>
	0xAD: [`\u833C`].string() // U+833C <cjk>
	0xAE: [`\u8344`].string() // U+8344 <cjk>
	0xAF: [`\u8357`].string() // U+8357 <cjk>
	0xB0: [`\u44BE`].string() // U+44BE <cjk>
	0xB1: [`\u837F`].string() // U+837F <cjk>
	0xB2: [`\u44D4`].string() // U+44D4 <cjk>
	0xB3: [`\u44B3`].string() // U+44B3 <cjk>
	0xB4: [`\u838D`].string() // U+838D <cjk>
	0xB5: [`\u8394`].string() // U+8394 <cjk>
	0xB6: [`\u8395`].string() // U+8395 <cjk>
	0xB7: [`\u839B`].string() // U+839B <cjk>
	0xB8: [`\u839D`].string() // U+839D <cjk>
	0xB9: [`\u83C9`].string() // U+83C9 <cjk>
	0xBA: [`\u83D0`].string() // U+83D0 <cjk>
	0xBB: [`\u83D4`].string() // U+83D4 <cjk>
	0xBC: [`\u83DD`].string() // U+83DD <cjk>
	0xBD: [`\u83E5`].string() // U+83E5 <cjk>
	0xBE: [`\u83F9`].string() // U+83F9 <cjk>
	0xBF: [`\u840F`].string() // U+840F <cjk>
	0xC0: [`\u8411`].string() // U+8411 <cjk>
	0xC1: [`\u8415`].string() // U+8415 <cjk>
	0xC2: utf32_to_str(0x26C73) // U+26C73 <cjk>
	0xC3: [`\u8417`].string() // U+8417 <cjk>
	0xC4: [`\u8439`].string() // U+8439 <cjk>
	0xC5: [`\u844A`].string() // U+844A <cjk>
	0xC6: [`\u844F`].string() // U+844F <cjk>
	0xC7: [`\u8451`].string() // U+8451 <cjk>
	0xC8: [`\u8452`].string() // U+8452 <cjk>
	0xC9: [`\u8459`].string() // U+8459 <cjk>
	0xCA: [`\u845A`].string() // U+845A <cjk>
	0xCB: [`\u845C`].string() // U+845C <cjk>
	0xCC: utf32_to_str(0x26CDD) // U+26CDD <cjk>
	0xCD: [`\u8465`].string() // U+8465 <cjk>
	0xCE: [`\u8476`].string() // U+8476 <cjk>
	0xCF: [`\u8478`].string() // U+8478 <cjk>
	0xD0: [`\u847C`].string() // U+847C <cjk>
	0xD1: [`\u8481`].string() // U+8481 <cjk>
	0xD2: [`\u450D`].string() // U+450D <cjk>
	0xD3: [`\u84DC`].string() // U+84DC <cjk>
	0xD4: [`\u8497`].string() // U+8497 <cjk>
	0xD5: [`\u84A6`].string() // U+84A6 <cjk>
	0xD6: [`\u84BE`].string() // U+84BE <cjk>
	0xD7: [`\u4508`].string() // U+4508 <cjk>
	0xD8: [`\u84CE`].string() // U+84CE <cjk>
	0xD9: [`\u84CF`].string() // U+84CF <cjk>
	0xDA: [`\u84D3`].string() // U+84D3 <cjk>
	0xDB: utf32_to_str(0x26E65) // U+26E65 <cjk>
	0xDC: [`\u84E7`].string() // U+84E7 <cjk>
	0xDD: [`\u84EA`].string() // U+84EA <cjk>
	0xDE: [`\u84EF`].string() // U+84EF <cjk>
	0xDF: [`\u84F0`].string() // U+84F0 <cjk>
	0xE0: [`\u84F1`].string() // U+84F1 <cjk>
	0xE1: [`\u84FA`].string() // U+84FA <cjk>
	0xE2: [`\u84FD`].string() // U+84FD <cjk>
	0xE3: [`\u850C`].string() // U+850C <cjk>
	0xE4: [`\u851B`].string() // U+851B <cjk>
	0xE5: [`\u8524`].string() // U+8524 <cjk>
	0xE6: [`\u8525`].string() // U+8525 <cjk>
	0xE7: [`\u852B`].string() // U+852B <cjk>
	0xE8: [`\u8534`].string() // U+8534 <cjk>
	0xE9: [`\u854F`].string() // U+854F <cjk>
	0xEA: [`\u856F`].string() // U+856F <cjk>
	0xEB: [`\u4525`].string() // U+4525 <cjk>
	0xEC: [`\u4543`].string() // U+4543 <cjk>
	0xED: [`\u853E`].string() // U+853E <cjk>
	0xEE: [`\u8551`].string() // U+8551 <cjk>
	0xEF: [`\u8553`].string() // U+8553 <cjk>
	0xF0: [`\u855E`].string() // U+855E <cjk>
	0xF1: [`\u8561`].string() // U+8561 <cjk>
	0xF2: [`\u8562`].string() // U+8562 <cjk>
	0xF3: utf32_to_str(0x26F94) // U+26F94 <cjk>
	0xF4: [`\u857B`].string() // U+857B <cjk>
	0xF5: [`\u857D`].string() // U+857D <cjk>
	0xF6: [`\u857F`].string() // U+857F <cjk>
	0xF7: [`\u8581`].string() // U+8581 <cjk>
	0xF8: [`\u8586`].string() // U+8586 <cjk>
	0xF9: [`\u8593`].string() // U+8593 <cjk>
	0xFA: [`\u859D`].string() // U+859D <cjk>
	0xFB: [`\u859F`].string() // U+859F <cjk>
	0xFC: utf32_to_str(0x26FF8) // U+26FF8 <cjk>
}

module mojibake

const jis_x_0213_doublebyte_0x8b = {
	0x40: [`\u6A5F`].string() // U+6A5F <cjk>
	0x41: [`\u5E30`].string() // U+5E30 <cjk>
	0x42: [`\u6BC5`].string() // U+6BC5 <cjk>
	0x43: [`\u6C17`].string() // U+6C17 <cjk>
	0x44: [`\u6C7D`].string() // U+6C7D <cjk>
	0x45: [`\u757F`].string() // U+757F <cjk>
	0x46: [`\u7948`].string() // U+7948 <cjk>
	0x47: [`\u5B63`].string() // U+5B63 <cjk>
	0x48: [`\u7A00`].string() // U+7A00 <cjk>
	0x49: [`\u7D00`].string() // U+7D00 <cjk>
	0x4A: [`\u5FBD`].string() // U+5FBD <cjk>
	0x4B: [`\u898F`].string() // U+898F <cjk>
	0x4C: [`\u8A18`].string() // U+8A18 <cjk>
	0x4D: [`\u8CB4`].string() // U+8CB4 <cjk>
	0x4E: [`\u8D77`].string() // U+8D77 <cjk>
	0x4F: [`\u8ECC`].string() // U+8ECC <cjk>
	0x50: [`\u8F1D`].string() // U+8F1D <cjk>
	0x51: [`\u98E2`].string() // U+98E2 <cjk>
	0x52: [`\u9A0E`].string() // U+9A0E <cjk>
	0x53: [`\u9B3C`].string() // U+9B3C <cjk>
	0x54: [`\u4E80`].string() // U+4E80 <cjk>
	0x55: [`\u507D`].string() // U+507D <cjk>
	0x56: [`\u5100`].string() // U+5100 <cjk>
	0x57: [`\u5993`].string() // U+5993 <cjk>
	0x58: [`\u5B9C`].string() // U+5B9C <cjk>
	0x59: [`\u622F`].string() // U+622F <cjk>
	0x5A: [`\u6280`].string() // U+6280 <cjk>
	0x5B: [`\u64EC`].string() // U+64EC <cjk>
	0x5C: [`\u6B3A`].string() // U+6B3A <cjk>
	0x5D: [`\u72A0`].string() // U+72A0 <cjk>
	0x5E: [`\u7591`].string() // U+7591 <cjk>
	0x5F: [`\u7947`].string() // U+7947 <cjk>
	0x60: [`\u7FA9`].string() // U+7FA9 <cjk>
	0x61: [`\u87FB`].string() // U+87FB <cjk>
	0x62: [`\u8ABC`].string() // U+8ABC <cjk>
	0x63: [`\u8B70`].string() // U+8B70 <cjk>
	0x64: [`\u63AC`].string() // U+63AC <cjk>
	0x65: [`\u83CA`].string() // U+83CA <cjk>
	0x66: [`\u97A0`].string() // U+97A0 <cjk>
	0x67: [`\u5409`].string() // U+5409 <cjk>
	0x68: [`\u5403`].string() // U+5403 <cjk>
	0x69: [`\u55AB`].string() // U+55AB <cjk>
	0x6A: [`\u6854`].string() // U+6854 <cjk>
	0x6B: [`\u6A58`].string() // U+6A58 <cjk>
	0x6C: [`\u8A70`].string() // U+8A70 <cjk>
	0x6D: [`\u7827`].string() // U+7827 <cjk>
	0x6E: [`\u6775`].string() // U+6775 <cjk>
	0x6F: [`\u9ECD`].string() // U+9ECD <cjk>
	0x70: [`\u5374`].string() // U+5374 <cjk>
	0x71: [`\u5BA2`].string() // U+5BA2 <cjk>
	0x72: [`\u811A`].string() // U+811A <cjk>
	0x73: [`\u8650`].string() // U+8650 <cjk>
	0x74: [`\u9006`].string() // U+9006 <cjk>
	0x75: [`\u4E18`].string() // U+4E18 <cjk>
	0x76: [`\u4E45`].string() // U+4E45 <cjk>
	0x77: [`\u4EC7`].string() // U+4EC7 <cjk>
	0x78: [`\u4F11`].string() // U+4F11 <cjk>
	0x79: [`\u53CA`].string() // U+53CA <cjk>
	0x7A: [`\u5438`].string() // U+5438 <cjk>
	0x7B: [`\u5BAE`].string() // U+5BAE <cjk>
	0x7C: [`\u5F13`].string() // U+5F13 <cjk>
	0x7D: [`\u6025`].string() // U+6025 <cjk>
	0x7E: [`\u6551`].string() // U+6551 <cjk>
	0x80: [`\u673D`].string() // U+673D <cjk>
	0x81: [`\u6C42`].string() // U+6C42 <cjk>
	0x82: [`\u6C72`].string() // U+6C72 <cjk>
	0x83: [`\u6CE3`].string() // U+6CE3 <cjk>
	0x84: [`\u7078`].string() // U+7078 <cjk>
	0x85: [`\u7403`].string() // U+7403 <cjk>
	0x86: [`\u7A76`].string() // U+7A76 <cjk>
	0x87: [`\u7AAE`].string() // U+7AAE <cjk>
	0x88: [`\u7B08`].string() // U+7B08 <cjk>
	0x89: [`\u7D1A`].string() // U+7D1A <cjk>
	0x8A: [`\u7CFE`].string() // U+7CFE <cjk>
	0x8B: [`\u7D66`].string() // U+7D66 <cjk>
	0x8C: [`\u65E7`].string() // U+65E7 <cjk>
	0x8D: [`\u725B`].string() // U+725B <cjk>
	0x8E: [`\u53BB`].string() // U+53BB <cjk>
	0x8F: [`\u5C45`].string() // U+5C45 <cjk>
	0x90: [`\u5DE8`].string() // U+5DE8 <cjk>
	0x91: [`\u62D2`].string() // U+62D2 <cjk>
	0x92: [`\u62E0`].string() // U+62E0 <cjk>
	0x93: [`\u6319`].string() // U+6319 <cjk>
	0x94: [`\u6E20`].string() // U+6E20 <cjk>
	0x95: [`\u865A`].string() // U+865A <cjk>
	0x96: [`\u8A31`].string() // U+8A31 <cjk>
	0x97: [`\u8DDD`].string() // U+8DDD <cjk>
	0x98: [`\u92F8`].string() // U+92F8 <cjk>
	0x99: [`\u6F01`].string() // U+6F01 <cjk>
	0x9A: [`\u79A6`].string() // U+79A6 <cjk>
	0x9B: [`\u9B5A`].string() // U+9B5A <cjk>
	0x9C: [`\u4EA8`].string() // U+4EA8 <cjk>
	0x9D: [`\u4EAB`].string() // U+4EAB <cjk>
	0x9E: [`\u4EAC`].string() // U+4EAC <cjk>
	0x9F: [`\u4F9B`].string() // U+4F9B <cjk>
	0xA0: [`\u4FA0`].string() // U+4FA0 <cjk>
	0xA1: [`\u50D1`].string() // U+50D1 <cjk>
	0xA2: [`\u5147`].string() // U+5147 <cjk>
	0xA3: [`\u7AF6`].string() // U+7AF6 <cjk>
	0xA4: [`\u5171`].string() // U+5171 <cjk>
	0xA5: [`\u51F6`].string() // U+51F6 <cjk>
	0xA6: [`\u5354`].string() // U+5354 <cjk>
	0xA7: [`\u5321`].string() // U+5321 <cjk>
	0xA8: [`\u537F`].string() // U+537F <cjk>
	0xA9: [`\u53EB`].string() // U+53EB <cjk>
	0xAA: [`\u55AC`].string() // U+55AC <cjk>
	0xAB: [`\u5883`].string() // U+5883 <cjk>
	0xAC: [`\u5CE1`].string() // U+5CE1 <cjk>
	0xAD: [`\u5F37`].string() // U+5F37 <cjk>
	0xAE: [`\u5F4A`].string() // U+5F4A <cjk>
	0xAF: [`\u602F`].string() // U+602F <cjk>
	0xB0: [`\u6050`].string() // U+6050 <cjk>
	0xB1: [`\u606D`].string() // U+606D <cjk>
	0xB2: [`\u631F`].string() // U+631F <cjk>
	0xB3: [`\u6559`].string() // U+6559 <cjk>
	0xB4: [`\u6A4B`].string() // U+6A4B <cjk>
	0xB5: [`\u6CC1`].string() // U+6CC1 <cjk>
	0xB6: [`\u72C2`].string() // U+72C2 <cjk>
	0xB7: [`\u72ED`].string() // U+72ED <cjk>
	0xB8: [`\u77EF`].string() // U+77EF <cjk>
	0xB9: [`\u80F8`].string() // U+80F8 <cjk>
	0xBA: [`\u8105`].string() // U+8105 <cjk>
	0xBB: [`\u8208`].string() // U+8208 <cjk>
	0xBC: [`\u854E`].string() // U+854E <cjk>
	0xBD: [`\u90F7`].string() // U+90F7 <cjk>
	0xBE: [`\u93E1`].string() // U+93E1 <cjk>
	0xBF: [`\u97FF`].string() // U+97FF <cjk>
	0xC0: [`\u9957`].string() // U+9957 <cjk>
	0xC1: [`\u9A5A`].string() // U+9A5A <cjk>
	0xC2: [`\u4EF0`].string() // U+4EF0 <cjk>
	0xC3: [`\u51DD`].string() // U+51DD <cjk>
	0xC4: [`\u5C2D`].string() // U+5C2D <cjk>
	0xC5: [`\u6681`].string() // U+6681 <cjk>
	0xC6: [`\u696D`].string() // U+696D <cjk>
	0xC7: [`\u5C40`].string() // U+5C40 <cjk>
	0xC8: [`\u66F2`].string() // U+66F2 <cjk>
	0xC9: [`\u6975`].string() // U+6975 <cjk>
	0xCA: [`\u7389`].string() // U+7389 <cjk>
	0xCB: [`\u6850`].string() // U+6850 <cjk>
	0xCC: [`\u7C81`].string() // U+7C81 <cjk>
	0xCD: [`\u50C5`].string() // U+50C5 <cjk>
	0xCE: [`\u52E4`].string() // U+52E4 <cjk>
	0xCF: [`\u5747`].string() // U+5747 <cjk>
	0xD0: [`\u5DFE`].string() // U+5DFE <cjk>
	0xD1: [`\u9326`].string() // U+9326 <cjk>
	0xD2: [`\u65A4`].string() // U+65A4 <cjk>
	0xD3: [`\u6B23`].string() // U+6B23 <cjk>
	0xD4: [`\u6B3D`].string() // U+6B3D <cjk>
	0xD5: [`\u7434`].string() // U+7434 <cjk>
	0xD6: [`\u7981`].string() // U+7981 <cjk>
	0xD7: [`\u79BD`].string() // U+79BD <cjk>
	0xD8: [`\u7B4B`].string() // U+7B4B <cjk>
	0xD9: [`\u7DCA`].string() // U+7DCA <cjk>
	0xDA: [`\u82B9`].string() // U+82B9 <cjk>
	0xDB: [`\u83CC`].string() // U+83CC <cjk>
	0xDC: [`\u887F`].string() // U+887F <cjk>
	0xDD: [`\u895F`].string() // U+895F <cjk>
	0xDE: [`\u8B39`].string() // U+8B39 <cjk>
	0xDF: [`\u8FD1`].string() // U+8FD1 <cjk>
	0xE0: [`\u91D1`].string() // U+91D1 <cjk>
	0xE1: [`\u541F`].string() // U+541F <cjk>
	0xE2: [`\u9280`].string() // U+9280 <cjk>
	0xE3: [`\u4E5D`].string() // U+4E5D <cjk>
	0xE4: [`\u5036`].string() // U+5036 <cjk>
	0xE5: [`\u53E5`].string() // U+53E5 <cjk>
	0xE6: [`\u533A`].string() // U+533A <cjk>
	0xE7: [`\u72D7`].string() // U+72D7 <cjk>
	0xE8: [`\u7396`].string() // U+7396 <cjk>
	0xE9: [`\u77E9`].string() // U+77E9 <cjk>
	0xEA: [`\u82E6`].string() // U+82E6 <cjk>
	0xEB: [`\u8EAF`].string() // U+8EAF <cjk>
	0xEC: [`\u99C6`].string() // U+99C6 <cjk>
	0xED: [`\u99C8`].string() // U+99C8 <cjk>
	0xEE: [`\u99D2`].string() // U+99D2 <cjk>
	0xEF: [`\u5177`].string() // U+5177 <cjk>
	0xF0: [`\u611A`].string() // U+611A <cjk>
	0xF1: [`\u865E`].string() // U+865E <cjk>
	0xF2: [`\u55B0`].string() // U+55B0 <cjk>
	0xF3: [`\u7A7A`].string() // U+7A7A <cjk>
	0xF4: [`\u5076`].string() // U+5076 <cjk>
	0xF5: [`\u5BD3`].string() // U+5BD3 <cjk>
	0xF6: [`\u9047`].string() // U+9047 <cjk>
	0xF7: [`\u9685`].string() // U+9685 <cjk>
	0xF8: [`\u4E32`].string() // U+4E32 <cjk>
	0xF9: [`\u6ADB`].string() // U+6ADB <cjk>
	0xFA: [`\u91E7`].string() // U+91E7 <cjk>
	0xFB: [`\u5C51`].string() // U+5C51 <cjk>
	0xFC: [`\u5C48`].string() // U+5C48 <cjk>
}

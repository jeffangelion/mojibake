module mojibake

const jis_x_0213_doublebyte_0x85 = {
	0x40: [`\u20AC`].string() // U+20AC EURO SIGN
	0x41: [`\u00A0`].string() // U+00A0 NO-BREAK SPACE
	0x42: [`\u00A1`].string() // U+00A1 INVERTED EXCLAMATION MARK
	0x43: [`\u00A4`].string() // U+00A4 CURRENCY SIGN
	0x44: [`\u00A6`].string() // U+00A6 BROKEN BAR
	0x45: [`\u00A9`].string() // U+00A9 COPYRIGHT SIGN
	0x46: [`\u00AA`].string() // U+00AA FEMININE ORDINAL INDICATOR
	0x47: [`\u00AB`].string() // U+00AB LEFT-POINTING DOUBLE ANGLE QUOTATION MARK
	0x48: [`\u00AD`].string() // U+00AD SOFT HYPHEN
	0x49: [`\u00AE`].string() // U+00AE REGISTERED SIGN
	0x4A: [`\u00AF`].string() // U+00AF MACRON
	0x4B: [`\u00B2`].string() // U+00B2 SUPERSCRIPT TWO
	0x4C: [`\u00B3`].string() // U+00B3 SUPERSCRIPT THREE
	0x4D: [`\u00B7`].string() // U+00B7 MIDDLE DOT
	0x4E: [`\u00B8`].string() // U+00B8 CEDILLA
	0x4F: [`\u00B9`].string() // U+00B9 SUPERSCRIPT ONE
	0x50: [`\u00BA`].string() // U+00BA MASCULINE ORDINAL INDICATOR
	0x51: [`\u00BB`].string() // U+00BB RIGHT-POINTING DOUBLE ANGLE QUOTATION MARK
	0x52: [`\u00BC`].string() // U+00BC VULGAR FRACTION ONE QUARTER
	0x53: [`\u00BD`].string() // U+00BD VULGAR FRACTION ONE HALF
	0x54: [`\u00BE`].string() // U+00BE VULGAR FRACTION THREE QUARTERS
	0x55: [`\u00BF`].string() // U+00BF INVERTED QUESTION MARK
	0x56: [`\u00C0`].string() // U+00C0 LATIN CAPITAL LETTER A WITH GRAVE
	0x57: [`\u00C1`].string() // U+00C1 LATIN CAPITAL LETTER A WITH ACUTE
	0x58: [`\u00C2`].string() // U+00C2 LATIN CAPITAL LETTER A WITH CIRCUMFLEX
	0x59: [`\u00C3`].string() // U+00C3 LATIN CAPITAL LETTER A WITH TILDE
	0x5A: [`\u00C4`].string() // U+00C4 LATIN CAPITAL LETTER A WITH DIAERESIS
	0x5B: [`\u00C5`].string() // U+00C5 LATIN CAPITAL LETTER A WITH RING ABOVE
	0x5C: [`\u00C6`].string() // U+00C6 LATIN CAPITAL LETTER AE
	0x5D: [`\u00C7`].string() // U+00C7 LATIN CAPITAL LETTER C WITH CEDILLA
	0x5E: [`\u00C8`].string() // U+00C8 LATIN CAPITAL LETTER E WITH GRAVE
	0x5F: [`\u00C9`].string() // U+00C9 LATIN CAPITAL LETTER E WITH ACUTE
	0x60: [`\u00CA`].string() // U+00CA LATIN CAPITAL LETTER E WITH CIRCUMFLEX
	0x61: [`\u00CB`].string() // U+00CB LATIN CAPITAL LETTER E WITH DIAERESIS
	0x62: [`\u00CC`].string() // U+00CC LATIN CAPITAL LETTER I WITH GRAVE
	0x63: [`\u00CD`].string() // U+00CD LATIN CAPITAL LETTER I WITH ACUTE
	0x64: [`\u00CE`].string() // U+00CE LATIN CAPITAL LETTER I WITH CIRCUMFLEX
	0x65: [`\u00CF`].string() // U+00CF LATIN CAPITAL LETTER I WITH DIAERESIS
	0x66: [`\u00D0`].string() // U+00D0 LATIN CAPITAL LETTER ETH
	0x67: [`\u00D1`].string() // U+00D1 LATIN CAPITAL LETTER N WITH TILDE
	0x68: [`\u00D2`].string() // U+00D2 LATIN CAPITAL LETTER O WITH GRAVE
	0x69: [`\u00D3`].string() // U+00D3 LATIN CAPITAL LETTER O WITH ACUTE
	0x6A: [`\u00D4`].string() // U+00D4 LATIN CAPITAL LETTER O WITH CIRCUMFLEX
	0x6B: [`\u00D5`].string() // U+00D5 LATIN CAPITAL LETTER O WITH TILDE
	0x6C: [`\u00D6`].string() // U+00D6 LATIN CAPITAL LETTER O WITH DIAERESIS
	0x6D: [`\u00D8`].string() // U+00D8 LATIN CAPITAL LETTER O WITH STROKE
	0x6E: [`\u00D9`].string() // U+00D9 LATIN CAPITAL LETTER U WITH GRAVE
	0x6F: [`\u00DA`].string() // U+00DA LATIN CAPITAL LETTER U WITH ACUTE
	0x70: [`\u00DB`].string() // U+00DB LATIN CAPITAL LETTER U WITH CIRCUMFLEX
	0x71: [`\u00DC`].string() // U+00DC LATIN CAPITAL LETTER U WITH DIAERESIS
	0x72: [`\u00DD`].string() // U+00DD LATIN CAPITAL LETTER Y WITH ACUTE
	0x73: [`\u00DE`].string() // U+00DE LATIN CAPITAL LETTER THORN
	0x74: [`\u00DF`].string() // U+00DF LATIN SMALL LETTER SHARP S
	0x75: [`\u00E0`].string() // U+00E0 LATIN SMALL LETTER A WITH GRAVE
	0x76: [`\u00E1`].string() // U+00E1 LATIN SMALL LETTER A WITH ACUTE
	0x77: [`\u00E2`].string() // U+00E2 LATIN SMALL LETTER A WITH CIRCUMFLEX
	0x78: [`\u00E3`].string() // U+00E3 LATIN SMALL LETTER A WITH TILDE
	0x79: [`\u00E4`].string() // U+00E4 LATIN SMALL LETTER A WITH DIAERESIS
	0x7A: [`\u00E5`].string() // U+00E5 LATIN SMALL LETTER A WITH RING ABOVE
	0x7B: [`\u00E6`].string() // U+00E6 LATIN SMALL LETTER AE
	0x7C: [`\u00E7`].string() // U+00E7 LATIN SMALL LETTER C WITH CEDILLA
	0x7D: [`\u00E8`].string() // U+00E8 LATIN SMALL LETTER E WITH GRAVE
	0x7E: [`\u00E9`].string() // U+00E9 LATIN SMALL LETTER E WITH ACUTE
	0x80: [`\u00EA`].string() // U+00EA LATIN SMALL LETTER E WITH CIRCUMFLEX
	0x81: [`\u00EB`].string() // U+00EB LATIN SMALL LETTER E WITH DIAERESIS
	0x82: [`\u00EC`].string() // U+00EC LATIN SMALL LETTER I WITH GRAVE
	0x83: [`\u00ED`].string() // U+00ED LATIN SMALL LETTER I WITH ACUTE
	0x84: [`\u00EE`].string() // U+00EE LATIN SMALL LETTER I WITH CIRCUMFLEX
	0x85: [`\u00EF`].string() // U+00EF LATIN SMALL LETTER I WITH DIAERESIS
	0x86: [`\u00F0`].string() // U+00F0 LATIN SMALL LETTER ETH
	0x87: [`\u00F1`].string() // U+00F1 LATIN SMALL LETTER N WITH TILDE
	0x88: [`\u00F2`].string() // U+00F2 LATIN SMALL LETTER O WITH GRAVE
	0x89: [`\u00F3`].string() // U+00F3 LATIN SMALL LETTER O WITH ACUTE
	0x8A: [`\u00F4`].string() // U+00F4 LATIN SMALL LETTER O WITH CIRCUMFLEX
	0x8B: [`\u00F5`].string() // U+00F5 LATIN SMALL LETTER O WITH TILDE
	0x8C: [`\u00F6`].string() // U+00F6 LATIN SMALL LETTER O WITH DIAERESIS
	0x8D: [`\u00F8`].string() // U+00F8 LATIN SMALL LETTER O WITH STROKE
	0x8E: [`\u00F9`].string() // U+00F9 LATIN SMALL LETTER U WITH GRAVE
	0x8F: [`\u00FA`].string() // U+00FA LATIN SMALL LETTER U WITH ACUTE
	0x90: [`\u00FB`].string() // U+00FB LATIN SMALL LETTER U WITH CIRCUMFLEX
	0x91: [`\u00FC`].string() // U+00FC LATIN SMALL LETTER U WITH DIAERESIS
	0x92: [`\u00FD`].string() // U+00FD LATIN SMALL LETTER Y WITH ACUTE
	0x93: [`\u00FE`].string() // U+00FE LATIN SMALL LETTER THORN
	0x94: [`\u00FF`].string() // U+00FF LATIN SMALL LETTER Y WITH DIAERESIS
	0x95: [`\u0100`].string() // U+0100 LATIN CAPITAL LETTER A WITH MACRON
	0x96: [`\u012A`].string() // U+012A LATIN CAPITAL LETTER I WITH MACRON
	0x97: [`\u016A`].string() // U+016A LATIN CAPITAL LETTER U WITH MACRON
	0x98: [`\u0112`].string() // U+0112 LATIN CAPITAL LETTER E WITH MACRON
	0x99: [`\u014C`].string() // U+014C LATIN CAPITAL LETTER O WITH MACRON
	0x9A: [`\u0101`].string() // U+0101 LATIN SMALL LETTER A WITH MACRON
	0x9B: [`\u012B`].string() // U+012B LATIN SMALL LETTER I WITH MACRON
	0x9C: [`\u016B`].string() // U+016B LATIN SMALL LETTER U WITH MACRON
	0x9D: [`\u0113`].string() // U+0113 LATIN SMALL LETTER E WITH MACRON
	0x9E: [`\u014D`].string() // U+014D LATIN SMALL LETTER O WITH MACRON
	0x9F: [`\u0104`].string() // U+0104 LATIN CAPITAL LETTER A WITH OGONEK
	0xA0: [`\u02D8`].string() // U+02D8 BREVE
	0xA1: [`\u0141`].string() // U+0141 LATIN CAPITAL LETTER L WITH STROKE
	0xA2: [`\u013D`].string() // U+013D LATIN CAPITAL LETTER L WITH CARON
	0xA3: [`\u015A`].string() // U+015A LATIN CAPITAL LETTER S WITH ACUTE
	0xA4: [`\u0160`].string() // U+0160 LATIN CAPITAL LETTER S WITH CARON
	0xA5: [`\u015E`].string() // U+015E LATIN CAPITAL LETTER S WITH CEDILLA
	0xA6: [`\u0164`].string() // U+0164 LATIN CAPITAL LETTER T WITH CARON
	0xA7: [`\u0179`].string() // U+0179 LATIN CAPITAL LETTER Z WITH ACUTE
	0xA8: [`\u017D`].string() // U+017D LATIN CAPITAL LETTER Z WITH CARON
	0xA9: [`\u017B`].string() // U+017B LATIN CAPITAL LETTER Z WITH DOT ABOVE
	0xAA: [`\u0105`].string() // U+0105 LATIN SMALL LETTER A WITH OGONEK
	0xAB: [`\u02DB`].string() // U+02DB OGONEK
	0xAC: [`\u0142`].string() // U+0142 LATIN SMALL LETTER L WITH STROKE
	0xAD: [`\u013E`].string() // U+013E LATIN SMALL LETTER L WITH CARON
	0xAE: [`\u015B`].string() // U+015B LATIN SMALL LETTER S WITH ACUTE
	0xAF: [`\u02C7`].string() // U+02C7 CARON
	0xB0: [`\u0161`].string() // U+0161 LATIN SMALL LETTER S WITH CARON
	0xB1: [`\u015F`].string() // U+015F LATIN SMALL LETTER S WITH CEDILLA
	0xB2: [`\u0165`].string() // U+0165 LATIN SMALL LETTER T WITH CARON
	0xB3: [`\u017A`].string() // U+017A LATIN SMALL LETTER Z WITH ACUTE
	0xB4: [`\u02DD`].string() // U+02DD DOUBLE ACUTE ACCENT
	0xB5: [`\u017E`].string() // U+017E LATIN SMALL LETTER Z WITH CARON
	0xB6: [`\u017C`].string() // U+017C LATIN SMALL LETTER Z WITH DOT ABOVE
	0xB7: [`\u0154`].string() // U+0154 LATIN CAPITAL LETTER R WITH ACUTE
	0xB8: [`\u0102`].string() // U+0102 LATIN CAPITAL LETTER A WITH BREVE
	0xB9: [`\u0139`].string() // U+0139 LATIN CAPITAL LETTER L WITH ACUTE
	0xBA: [`\u0106`].string() // U+0106 LATIN CAPITAL LETTER C WITH ACUTE
	0xBB: [`\u010C`].string() // U+010C LATIN CAPITAL LETTER C WITH CARON
	0xBC: [`\u0118`].string() // U+0118 LATIN CAPITAL LETTER E WITH OGONEK
	0xBD: [`\u011A`].string() // U+011A LATIN CAPITAL LETTER E WITH CARON
	0xBE: [`\u010E`].string() // U+010E LATIN CAPITAL LETTER D WITH CARON
	0xBF: [`\u0143`].string() // U+0143 LATIN CAPITAL LETTER N WITH ACUTE
	0xC0: [`\u0147`].string() // U+0147 LATIN CAPITAL LETTER N WITH CARON
	0xC1: [`\u0150`].string() // U+0150 LATIN CAPITAL LETTER O WITH DOUBLE ACUTE
	0xC2: [`\u0158`].string() // U+0158 LATIN CAPITAL LETTER R WITH CARON
	0xC3: [`\u016E`].string() // U+016E LATIN CAPITAL LETTER U WITH RING ABOVE
	0xC4: [`\u0170`].string() // U+0170 LATIN CAPITAL LETTER U WITH DOUBLE ACUTE
	0xC5: [`\u0162`].string() // U+0162 LATIN CAPITAL LETTER T WITH CEDILLA
	0xC6: [`\u0155`].string() // U+0155 LATIN SMALL LETTER R WITH ACUTE
	0xC7: [`\u0103`].string() // U+0103 LATIN SMALL LETTER A WITH BREVE
	0xC8: [`\u013A`].string() // U+013A LATIN SMALL LETTER L WITH ACUTE
	0xC9: [`\u0107`].string() // U+0107 LATIN SMALL LETTER C WITH ACUTE
	0xCA: [`\u010D`].string() // U+010D LATIN SMALL LETTER C WITH CARON
	0xCB: [`\u0119`].string() // U+0119 LATIN SMALL LETTER E WITH OGONEK
	0xCC: [`\u011B`].string() // U+011B LATIN SMALL LETTER E WITH CARON
	0xCD: [`\u010F`].string() // U+010F LATIN SMALL LETTER D WITH CARON
	0xCE: [`\u0111`].string() // U+0111 LATIN SMALL LETTER D WITH STROKE
	0xCF: [`\u0144`].string() // U+0144 LATIN SMALL LETTER N WITH ACUTE
	0xD0: [`\u0148`].string() // U+0148 LATIN SMALL LETTER N WITH CARON
	0xD1: [`\u0151`].string() // U+0151 LATIN SMALL LETTER O WITH DOUBLE ACUTE
	0xD2: [`\u0159`].string() // U+0159 LATIN SMALL LETTER R WITH CARON
	0xD3: [`\u016F`].string() // U+016F LATIN SMALL LETTER U WITH RING ABOVE
	0xD4: [`\u0171`].string() // U+0171 LATIN SMALL LETTER U WITH DOUBLE ACUTE
	0xD5: [`\u0163`].string() // U+0163 LATIN SMALL LETTER T WITH CEDILLA
	0xD6: [`\u02D9`].string() // U+02D9 DOT ABOVE
	0xD7: [`\u0108`].string() // U+0108 LATIN CAPITAL LETTER C WITH CIRCUMFLEX
	0xD8: [`\u011C`].string() // U+011C LATIN CAPITAL LETTER G WITH CIRCUMFLEX
	0xD9: [`\u0124`].string() // U+0124 LATIN CAPITAL LETTER H WITH CIRCUMFLEX
	0xDA: [`\u0134`].string() // U+0134 LATIN CAPITAL LETTER J WITH CIRCUMFLEX
	0xDB: [`\u015C`].string() // U+015C LATIN CAPITAL LETTER S WITH CIRCUMFLEX
	0xDC: [`\u016C`].string() // U+016C LATIN CAPITAL LETTER U WITH BREVE
	0xDD: [`\u0109`].string() // U+0109 LATIN SMALL LETTER C WITH CIRCUMFLEX
	0xDE: [`\u011D`].string() // U+011D LATIN SMALL LETTER G WITH CIRCUMFLEX
	0xDF: [`\u0125`].string() // U+0125 LATIN SMALL LETTER H WITH CIRCUMFLEX
	0xE0: [`\u0135`].string() // U+0135 LATIN SMALL LETTER J WITH CIRCUMFLEX
	0xE1: [`\u015D`].string() // U+015D LATIN SMALL LETTER S WITH CIRCUMFLEX
	0xE2: [`\u016D`].string() // U+016D LATIN SMALL LETTER U WITH BREVE
	0xE3: [`\u0271`].string() // U+0271 LATIN SMALL LETTER M WITH HOOK
	0xE4: [`\u028B`].string() // U+028B LATIN SMALL LETTER V WITH HOOK
	0xE5: [`\u027E`].string() // U+027E LATIN SMALL LETTER R WITH FISHHOOK
	0xE6: [`\u0283`].string() // U+0283 LATIN SMALL LETTER ESH
	0xE7: [`\u0292`].string() // U+0292 LATIN SMALL LETTER EZH
	0xE8: [`\u026C`].string() // U+026C LATIN SMALL LETTER L WITH BELT
	0xE9: [`\u026E`].string() // U+026E LATIN SMALL LETTER LEZH
	0xEA: [`\u0279`].string() // U+0279 LATIN SMALL LETTER TURNED R
	0xEB: [`\u0288`].string() // U+0288 LATIN SMALL LETTER T WITH RETROFLEX HOOK
	0xEC: [`\u0256`].string() // U+0256 LATIN SMALL LETTER D WITH TAIL
	0xED: [`\u0273`].string() // U+0273 LATIN SMALL LETTER N WITH RETROFLEX HOOK
	0xEE: [`\u027D`].string() // U+027D LATIN SMALL LETTER R WITH TAIL
	0xEF: [`\u0282`].string() // U+0282 LATIN SMALL LETTER S WITH HOOK
	0xF0: [`\u0290`].string() // U+0290 LATIN SMALL LETTER Z WITH RETROFLEX HOOK
	0xF1: [`\u027B`].string() // U+027B LATIN SMALL LETTER TURNED R WITH HOOK
	0xF2: [`\u026D`].string() // U+026D LATIN SMALL LETTER L WITH RETROFLEX HOOK
	0xF3: [`\u025F`].string() // U+025F LATIN SMALL LETTER DOTLESS J WITH STROKE
	0xF4: [`\u0272`].string() // U+0272 LATIN SMALL LETTER N WITH LEFT HOOK
	0xF5: [`\u029D`].string() // U+029D LATIN SMALL LETTER J WITH CROSSED-TAIL
	0xF6: [`\u028E`].string() // U+028E LATIN SMALL LETTER TURNED Y
	0xF7: [`\u0261`].string() // U+0261 LATIN SMALL LETTER SCRIPT G
	0xF8: [`\u014B`].string() // U+014B LATIN SMALL LETTER ENG
	0xF9: [`\u0270`].string() // U+0270 LATIN SMALL LETTER TURNED M WITH LONG LEG
	0xFA: [`\u0281`].string() // U+0281 LATIN LETTER SMALL CAPITAL INVERTED R
	0xFB: [`\u0127`].string() // U+0127 LATIN SMALL LETTER H WITH STROKE
	0xFC: [`\u0295`].string() // U+0295 LATIN LETTER PHARYNGEAL VOICED FRICATIVE
}
